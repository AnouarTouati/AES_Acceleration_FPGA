// ============================================================================

`define ENABLE_HPS
//`define ENABLE_HSMC

module DE10_Standard_GHRD(


      ///////// CLOCK /////////
      input              CLOCK2_50,
      input              CLOCK3_50,
      input              CLOCK4_50,
      input              CLOCK_50,

      ///////// KEY /////////
      input    [ 3: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LED /////////
      output   [ 9: 0]   LEDR,

      ///////// Seg7 /////////
      output   [ 6: 0]   HEX0,
      output   [ 6: 0]   HEX1,
      output   [ 6: 0]   HEX2,
      output   [ 6: 0]   HEX3,
      output   [ 6: 0]   HEX4,
      output   [ 6: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// Video-In /////////
      input              TD_CLK27,
      input              TD_HS,
      input              TD_VS,
      input    [ 7: 0]   TD_DATA,
      output             TD_RESET_N,

      ///////// VGA /////////
      output             VGA_CLK,
      output             VGA_HS,
      output             VGA_VS,
      output   [ 7: 0]   VGA_R,
      output   [ 7: 0]   VGA_G,
      output   [ 7: 0]   VGA_B,
      output             VGA_BLANK_N,
      output             VGA_SYNC_N,

      ///////// Audio /////////
      inout              AUD_BCLK,
      output             AUD_XCK,
      inout              AUD_ADCLRCK,
      input              AUD_ADCDAT,
      inout              AUD_DACLRCK,
      output             AUD_DACDAT,

      ///////// PS2 /////////
      inout              PS2_CLK,
      inout              PS2_CLK2,
      inout              PS2_DAT,
      inout              PS2_DAT2,

      ///////// ADC /////////
      output             ADC_SCLK,
      input              ADC_DOUT,
      output             ADC_DIN,
      output             ADC_CONVST,

      ///////// I2C for Audio and Video-In /////////
      output             FPGA_I2C_SCLK,
      inout              FPGA_I2C_SDAT,

      ///////// GPIO /////////
      inout    [35: 0]   GPIO,

`ifdef ENABLE_HSMC
      ///////// HSMC /////////
      input              HSMC_CLKIN_P1,
      input              HSMC_CLKIN_N1,
      input              HSMC_CLKIN_P2,
      input              HSMC_CLKIN_N2,
      output             HSMC_CLKOUT_P1,
      output             HSMC_CLKOUT_N1,
      output             HSMC_CLKOUT_P2,
      output             HSMC_CLKOUT_N2,
      inout    [16: 0]   HSMC_TX_D_P,
      inout    [16: 0]   HSMC_TX_D_N,
      inout    [16: 0]   HSMC_RX_D_P,
      inout    [16: 0]   HSMC_RX_D_N,
      input              HSMC_CLKIN0,
      output             HSMC_CLKOUT0,
      inout    [ 3: 0]   HSMC_D,
      output             HSMC_SCL,
      inout              HSMC_SDA,
`endif /*ENABLE_HSMC*/

`ifdef ENABLE_HPS
      ///////// HPS /////////
      inout              HPS_CONV_USB_N,
      output      [14:0] HPS_DDR3_ADDR,
      output      [2:0]  HPS_DDR3_BA,
      output             HPS_DDR3_CAS_N,
      output             HPS_DDR3_CKE,
      output             HPS_DDR3_CK_N,
      output             HPS_DDR3_CK_P,
      output             HPS_DDR3_CS_N,
      output      [3:0]  HPS_DDR3_DM,
      inout       [31:0] HPS_DDR3_DQ,
      inout       [3:0]  HPS_DDR3_DQS_N,
      inout       [3:0]  HPS_DDR3_DQS_P,
      output             HPS_DDR3_ODT,
      output             HPS_DDR3_RAS_N,
      output             HPS_DDR3_RESET_N,
      input              HPS_DDR3_RZQ,
      output             HPS_DDR3_WE_N,
      output             HPS_ENET_GTX_CLK,
      inout              HPS_ENET_INT_N,
      output             HPS_ENET_MDC,
      inout              HPS_ENET_MDIO,
      input              HPS_ENET_RX_CLK,
      input       [3:0]  HPS_ENET_RX_DATA,
      input              HPS_ENET_RX_DV,
      output      [3:0]  HPS_ENET_TX_DATA,
      output             HPS_ENET_TX_EN,
      inout       [3:0]  HPS_FLASH_DATA,
      output             HPS_FLASH_DCLK,
      output             HPS_FLASH_NCSO,
      inout              HPS_GSENSOR_INT,
      inout              HPS_I2C1_SCLK,
      inout              HPS_I2C1_SDAT,
      inout              HPS_I2C2_SCLK,
      inout              HPS_I2C2_SDAT,
      inout              HPS_I2C_CONTROL,
      inout              HPS_KEY,
      inout              HPS_LCM_BK,
      inout              HPS_LCM_D_C,
      inout              HPS_LCM_RST_N,
      output             HPS_LCM_SPIM_CLK,
      output             HPS_LCM_SPIM_MOSI,
      output             HPS_LCM_SPIM_SS,
		input 				 HPS_LCM_SPIM_MISO,
      inout              HPS_LED,
      inout              HPS_LTC_GPIO,
      output             HPS_SD_CLK,
      inout              HPS_SD_CMD,
      inout       [3:0]  HPS_SD_DATA,
      output             HPS_SPIM_CLK,
      input              HPS_SPIM_MISO,
      output             HPS_SPIM_MOSI,
      inout              HPS_SPIM_SS,
      input              HPS_UART_RX,
      output             HPS_UART_TX,
      input              HPS_USB_CLKOUT,
      inout       [7:0]  HPS_USB_DATA,
      input              HPS_USB_DIR,
      input              HPS_USB_NXT,
      output             HPS_USB_STP,
`endif /*ENABLE_HPS*/
      ///////// IR /////////
      output             IRDA_TXD,
      input              IRDA_RXD
);



//=======================================================
//  REG/WIRE declarations
//=======================================================
  wire  			hps_fpga_reset_n;
  wire [3:0] 	fpga_debounced_buttons;
  wire [8:0]  	fpga_led_internal;
  wire [2:0]  	hps_reset_req;
  wire        	hps_cold_reset;
  wire        	hps_warm_reset;
  wire        	hps_debug_reset;
  wire [27:0] 	stm_hw_events;
  wire        	fpga_clk_50;
  
  //interface module
//  wire [127:0] read_bus;
//  wire [127:0] write_bus;
//  wire [5:0]   addr_bus;
//  wire         write_s;
//  wire         read_s;
//  wire         ackn_s;
//  wire [15:0]  byte_en;
  
//  //aes core
//  wire [3:0]   control;//bit3: start -- bit2: load -- bit1: mode -- bit0: reset
//  wire [127:0] key_aes_core;
//  wire [127:0] data_in_aes_core;
//  wire [127:0] data_out_aes_core;
//  wire 			done;

  //pll
 // wire 				 pll_clk;
   
  
// connection of internal logics
  //assign LEDR[9:1] = fpga_led_internal;
  assign stm_hw_events    = {{4{1'b0}}, SW, fpga_led_internal, fpga_debounced_buttons};
  assign fpga_clk_50=CLOCK_50;
  
//=======================================================
wire   locked;
// vga
wire       vga_clk;
wire       vga_hs;
wire       vga_vs;
wire [7:0] vga_r;
wire [7:0] vga_g;
wire [7:0] vga_b;
//	For Audio CODEC
wire		AUD_CTRL_CLK;	//	For Audio Controller		
// vga on board
assign {VGA_R, VGA_G, VGA_B} = {vga_r,vga_g,vga_b};
assign VGA_BLANK_N = 1'b1;
assign VGA_SYNC_N = 1'b0;
assign VGA_HS = ~vga_hs;
assign VGA_VS = ~vga_vs;
assign VGA_CLK = vga_clk;
//=======================================================
  
  
//=======================================================
//  Structural coding
//=======================================================

//aes128_fast u1(
//      .clk      (pll_clk), 
//      .reset    (control[0]), 
//      .start    (control[3]), 
//      .mode     (control[1]), 
//      .load     (control[2]), 
//      .key      (key_aes_core), 
//      .data_in  (data_in_aes_core), 
//      .data_out (data_out_aes_core), 
//      .done     (done)
//);

//interfacing_module u2 (
//.clk             (pll_clk),
//.read_data_bus   (read_bus),
//.write_data_bus  (write_bus),
//.addr_data_bus   (addr_bus),
//.write_signal    (write_s),
//.byteenable		  (byte_en),
//.read_signal     (read_s),
//.ackn_signal     (ackn_s),
//
//
//.reset_aes       (reset_aes_core),
//.start_aes       (start_aes_core),
//.mode_aes        (mode_aes_core),
//.load_aes        (load_aes_core),
//.key_aes         (key_aes_core),
//.data_in_aes     (data_in_aes_core),
//.data_out_aes    (data_out_aes_core),
//.done_aes        (done_aes_core)
//);

soc_system u0 (      
		  .clk_clk                               (CLOCK_50),                             //                clk.clk
		  .reset_reset_n                         (1'b1),                                 //                reset.reset_n
		 
		 //clocks
		/*output wire  */   // .clk_sdram_clk(DRAM_CLK), 
		/*output wire  */   // .clk_vga_clk(vga_clk), 
		/*output wire  */   // .clk_aud_clk(AUD_CTRL_CLK), 
		//.audio_and_video_config_0_external_interface_SDAT  (FPGA_I2C_SDAT),        // audio_and_video_config_0_external_interface.SDAT
     // .audio_and_video_config_0_external_interface_SCLK   (FPGA_I2C_SCLK),    
		
// sdram buffer
		/*output wire [12:0] */    //.sdram_wire_addr(DRAM_ADDR),                                 
		/*output wire [1:0]  */    //.sdram_wire_ba(DRAM_BA),                                   
		/*output wire        */    //.sdram_wire_cas_n(DRAM_CAS_N),                                
		/*output wire        */    //.sdram_wire_cke(DRAM_CKE),                                  
		/*output wire        */    //.sdram_wire_cs_n(DRAM_CS_N),                                 
		/*inout  wire [15:0] */    //.sdram_wire_dq(DRAM_DQ),                                   
		/*output wire [1:0]  */    //.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),                                  
		/*output wire        */    //.sdram_wire_ras_n(DRAM_RAS_N),                                
		/*output wire        */    //.sdram_wire_we_n(DRAM_WE_N),    

	//TV in
      /*input  wire        */    //.alt_vip_cl_cvi_0_clocked_video_vid_clk(TD_CLK27),            
		/*input  wire [7:0]  */    //.alt_vip_cl_cvi_0_clocked_video_vid_data(TD_DATA),           
		/*input  wire        */    //.alt_vip_cl_cvi_0_clocked_video_vid_de(1'b1),             
		/*input  wire        */    //.alt_vip_cl_cvi_0_clocked_video_vid_datavalid(1'b1),      
		/*input  wire        */    //.alt_vip_cl_cvi_0_clocked_video_vid_locked(1'b1),         
		/*input  wire        */    //.alt_vip_cl_cvi_0_clocked_video_vid_f(),              
		/*input  wire        */    //.alt_vip_cl_cvi_0_clocked_video_vid_v_sync(),         
		/*input  wire        */    //.alt_vip_cl_cvi_0_clocked_video_vid_h_sync(),         
		/*input  wire [7:0]  */    //.alt_vip_cl_cvi_0_clocked_video_vid_color_encoding(), 
		/*input  wire [7:0]  */    //.alt_vip_cl_cvi_0_clocked_video_vid_bit_width(),      
		/*output wire        */    //.alt_vip_cl_cvi_0_clocked_video_sof(),                
		/*output wire        */    //.alt_vip_cl_cvi_0_clocked_video_sof_locked(),         
		/*output wire        */    //.alt_vip_cl_cvi_0_clocked_video_refclk_div(),         
		/*output wire        */    //.alt_vip_cl_cvi_0_clocked_video_clipping(),           
		/*output wire        */    //.alt_vip_cl_cvi_0_clocked_video_padding(),            
		/*output wire        */    //.alt_vip_cl_cvi_0_clocked_video_overflow(),        


		  //HPS ddr3
		  .memory_mem_a                          ( HPS_DDR3_ADDR),                       //                memory.mem_a
        .memory_mem_ba                         ( HPS_DDR3_BA),                         //                .mem_ba
        .memory_mem_ck                         ( HPS_DDR3_CK_P),                       //                .mem_ck
        .memory_mem_ck_n                       ( HPS_DDR3_CK_N),                       //                .mem_ck_n
        .memory_mem_cke                        ( HPS_DDR3_CKE),                        //                .mem_cke
        .memory_mem_cs_n                       ( HPS_DDR3_CS_N),                       //                .mem_cs_n
        .memory_mem_ras_n                      ( HPS_DDR3_RAS_N),                      //                .mem_ras_n
        .memory_mem_cas_n                      ( HPS_DDR3_CAS_N),                      //                .mem_cas_n
        .memory_mem_we_n                       ( HPS_DDR3_WE_N),                       //                .mem_we_n
        .memory_mem_reset_n                    ( HPS_DDR3_RESET_N),                    //                .mem_reset_n
        .memory_mem_dq                         ( HPS_DDR3_DQ),                         //                .mem_dq
        .memory_mem_dqs                        ( HPS_DDR3_DQS_P),                      //                .mem_dqs
        .memory_mem_dqs_n                      ( HPS_DDR3_DQS_N),                      //                .mem_dqs_n
        .memory_mem_odt                        ( HPS_DDR3_ODT),                        //                .mem_odt
        .memory_mem_dm                         ( HPS_DDR3_DM),                         //                .mem_dm
        .memory_oct_rzqin                      ( HPS_DDR3_RZQ),                        //                .oct_rzqin
       //HPS ethernet		
	     .hps_0_hps_io_hps_io_emac1_inst_TX_CLK ( HPS_ENET_GTX_CLK),       //                             hps_0_hps_io.hps_io_emac1_inst_TX_CLK
        .hps_0_hps_io_hps_io_emac1_inst_TXD0   ( HPS_ENET_TX_DATA[0] ),   //                             .hps_io_emac1_inst_TXD0
        .hps_0_hps_io_hps_io_emac1_inst_TXD1   ( HPS_ENET_TX_DATA[1] ),   //                             .hps_io_emac1_inst_TXD1
        .hps_0_hps_io_hps_io_emac1_inst_TXD2   ( HPS_ENET_TX_DATA[2] ),   //                             .hps_io_emac1_inst_TXD2
        .hps_0_hps_io_hps_io_emac1_inst_TXD3   ( HPS_ENET_TX_DATA[3] ),   //                             .hps_io_emac1_inst_TXD3
        .hps_0_hps_io_hps_io_emac1_inst_RXD0   ( HPS_ENET_RX_DATA[0] ),   //                             .hps_io_emac1_inst_RXD0
        .hps_0_hps_io_hps_io_emac1_inst_MDIO   ( HPS_ENET_MDIO ),         //                             .hps_io_emac1_inst_MDIO
        .hps_0_hps_io_hps_io_emac1_inst_MDC    ( HPS_ENET_MDC  ),         //                             .hps_io_emac1_inst_MDC
        .hps_0_hps_io_hps_io_emac1_inst_RX_CTL ( HPS_ENET_RX_DV),         //                             .hps_io_emac1_inst_RX_CTL
        .hps_0_hps_io_hps_io_emac1_inst_TX_CTL ( HPS_ENET_TX_EN),         //                             .hps_io_emac1_inst_TX_CTL
        .hps_0_hps_io_hps_io_emac1_inst_RX_CLK ( HPS_ENET_RX_CLK),        //                             .hps_io_emac1_inst_RX_CLK
        .hps_0_hps_io_hps_io_emac1_inst_RXD1   ( HPS_ENET_RX_DATA[1] ),   //                             .hps_io_emac1_inst_RXD1
        .hps_0_hps_io_hps_io_emac1_inst_RXD2   ( HPS_ENET_RX_DATA[2] ),   //                             .hps_io_emac1_inst_RXD2
        .hps_0_hps_io_hps_io_emac1_inst_RXD3   ( HPS_ENET_RX_DATA[3] ),   //                             .hps_io_emac1_inst_RXD3
       //HPS QSPI  
		  .hps_0_hps_io_hps_io_qspi_inst_IO0     ( HPS_FLASH_DATA[0]    ),     //                               .hps_io_qspi_inst_IO0
        .hps_0_hps_io_hps_io_qspi_inst_IO1     ( HPS_FLASH_DATA[1]    ),     //                               .hps_io_qspi_inst_IO1
        .hps_0_hps_io_hps_io_qspi_inst_IO2     ( HPS_FLASH_DATA[2]    ),     //                               .hps_io_qspi_inst_IO2
        .hps_0_hps_io_hps_io_qspi_inst_IO3     ( HPS_FLASH_DATA[3]    ),     //                               .hps_io_qspi_inst_IO3
        .hps_0_hps_io_hps_io_qspi_inst_SS0     ( HPS_FLASH_NCSO    ),        //                               .hps_io_qspi_inst_SS0
        .hps_0_hps_io_hps_io_qspi_inst_CLK     ( HPS_FLASH_DCLK    ),        //                               .hps_io_qspi_inst_CLK
       //HPS SD card 
		  .hps_0_hps_io_hps_io_sdio_inst_CMD     ( HPS_SD_CMD    ),           //                               .hps_io_sdio_inst_CMD
        .hps_0_hps_io_hps_io_sdio_inst_D0      ( HPS_SD_DATA[0]     ),      //                               .hps_io_sdio_inst_D0
        .hps_0_hps_io_hps_io_sdio_inst_D1      ( HPS_SD_DATA[1]     ),      //                               .hps_io_sdio_inst_D1
        .hps_0_hps_io_hps_io_sdio_inst_CLK     ( HPS_SD_CLK   ),            //                               .hps_io_sdio_inst_CLK
        .hps_0_hps_io_hps_io_sdio_inst_D2      ( HPS_SD_DATA[2]     ),      //                               .hps_io_sdio_inst_D2
        .hps_0_hps_io_hps_io_sdio_inst_D3      ( HPS_SD_DATA[3]     ),      //                               .hps_io_sdio_inst_D3
       //HPS USB 		  
		  .hps_0_hps_io_hps_io_usb1_inst_D0      ( HPS_USB_DATA[0]    ),      //                               .hps_io_usb1_inst_D0
        .hps_0_hps_io_hps_io_usb1_inst_D1      ( HPS_USB_DATA[1]    ),      //                               .hps_io_usb1_inst_D1
        .hps_0_hps_io_hps_io_usb1_inst_D2      ( HPS_USB_DATA[2]    ),      //                               .hps_io_usb1_inst_D2
        .hps_0_hps_io_hps_io_usb1_inst_D3      ( HPS_USB_DATA[3]    ),      //                               .hps_io_usb1_inst_D3
        .hps_0_hps_io_hps_io_usb1_inst_D4      ( HPS_USB_DATA[4]    ),      //                               .hps_io_usb1_inst_D4
        .hps_0_hps_io_hps_io_usb1_inst_D5      ( HPS_USB_DATA[5]    ),      //                               .hps_io_usb1_inst_D5
        .hps_0_hps_io_hps_io_usb1_inst_D6      ( HPS_USB_DATA[6]    ),      //                               .hps_io_usb1_inst_D6
        .hps_0_hps_io_hps_io_usb1_inst_D7      ( HPS_USB_DATA[7]    ),      //                               .hps_io_usb1_inst_D7
        .hps_0_hps_io_hps_io_usb1_inst_CLK     ( HPS_USB_CLKOUT    ),       //                               .hps_io_usb1_inst_CLK
        .hps_0_hps_io_hps_io_usb1_inst_STP     ( HPS_USB_STP    ),          //                               .hps_io_usb1_inst_STP
        .hps_0_hps_io_hps_io_usb1_inst_DIR     ( HPS_USB_DIR    ),          //                               .hps_io_usb1_inst_DIR
        .hps_0_hps_io_hps_io_usb1_inst_NXT     ( HPS_USB_NXT    ),          //                               .hps_io_usb1_inst_NXT
		  
		  //HPS SPI0->LCDM 	
        .hps_0_hps_io_hps_io_spim0_inst_CLK    ( HPS_LCM_SPIM_CLK),    //                               .hps_io_spim0_inst_CLK
        .hps_0_hps_io_hps_io_spim0_inst_MOSI   ( HPS_LCM_SPIM_MOSI),   //                               .hps_io_spim0_inst_MOSI
        .hps_0_hps_io_hps_io_spim0_inst_MISO   ( HPS_LCM_SPIM_MISO),   //                               .hps_io_spim0_inst_MISO
        .hps_0_hps_io_hps_io_spim0_inst_SS0    ( HPS_LCM_SPIM_SS),    //                               .hps_io_spim0_inst_SS0
       //HPS SPI1 		  
		  .hps_0_hps_io_hps_io_spim1_inst_CLK    ( HPS_SPIM_CLK  ),           //                               .hps_io_spim1_inst_CLK
        .hps_0_hps_io_hps_io_spim1_inst_MOSI   ( HPS_SPIM_MOSI ),           //                               .hps_io_spim1_inst_MOSI
        .hps_0_hps_io_hps_io_spim1_inst_MISO   ( HPS_SPIM_MISO ),           //                               .hps_io_spim1_inst_MISO
        .hps_0_hps_io_hps_io_spim1_inst_SS0    ( HPS_SPIM_SS ),             //                               .hps_io_spim1_inst_SS0
      //HPS UART		
		  .hps_0_hps_io_hps_io_uart0_inst_RX     ( HPS_UART_RX    ),          //                               .hps_io_uart0_inst_RX
        .hps_0_hps_io_hps_io_uart0_inst_TX     ( HPS_UART_TX    ),          //                               .hps_io_uart0_inst_TX
		//HPS I2C1
		  .hps_0_hps_io_hps_io_i2c0_inst_SDA     ( HPS_I2C1_SDAT    ),        //                               .hps_io_i2c0_inst_SDA
        .hps_0_hps_io_hps_io_i2c0_inst_SCL     ( HPS_I2C1_SCLK    ),        //                               .hps_io_i2c0_inst_SCL
		//HPS I2C2
		  .hps_0_hps_io_hps_io_i2c1_inst_SDA     ( HPS_I2C2_SDAT    ),        //                               .hps_io_i2c1_inst_SDA
        .hps_0_hps_io_hps_io_i2c1_inst_SCL     ( HPS_I2C2_SCLK    ),        //                               .hps_io_i2c1_inst_SCL
      //HPS GPIO  
		  .hps_0_hps_io_hps_io_gpio_inst_GPIO09  ( HPS_CONV_USB_N),           //                               .hps_io_gpio_inst_GPIO09
        .hps_0_hps_io_hps_io_gpio_inst_GPIO35  ( HPS_ENET_INT_N),           //                               .hps_io_gpio_inst_GPIO35
        .hps_0_hps_io_hps_io_gpio_inst_GPIO37  ( HPS_LCM_BK ),  //                               .hps_io_gpio_inst_GPIO37
		  .hps_0_hps_io_hps_io_gpio_inst_GPIO40  ( HPS_LTC_GPIO ),              //                               .hps_io_gpio_inst_GPIO40
        .hps_0_hps_io_hps_io_gpio_inst_GPIO41  ( HPS_LCM_D_C ),              //                               .hps_io_gpio_inst_GPIO41
        .hps_0_hps_io_hps_io_gpio_inst_GPIO44  ( HPS_LCM_RST_N  ),  //                               .hps_io_gpio_inst_GPIO44
		  .hps_0_hps_io_hps_io_gpio_inst_GPIO48  ( HPS_I2C_CONTROL),          //                               .hps_io_gpio_inst_GPIO48
        .hps_0_hps_io_hps_io_gpio_inst_GPIO53  ( HPS_LED),                  //                               .hps_io_gpio_inst_GPIO53
        .hps_0_hps_io_hps_io_gpio_inst_GPIO54  ( HPS_KEY),                  //                               .hps_io_gpio_inst_GPIO54
    	  .hps_0_hps_io_hps_io_gpio_inst_GPIO61  ( HPS_GSENSOR_INT),  //                               .hps_io_gpio_inst_GPIO61

			
		  //.led_pio_external_connection_export    ( fpga_led_internal ),               //                               led_pio_external_connection.export                     
        .dipsw_pio_external_connection_export  ( SW ),                 //                               dipsw_pio_external_connection.export
        .button_pio_external_connection_export ( fpga_debounced_buttons ),              //                               button_pio_external_connection.export 
		  //.hps_0_h2f_reset_reset_n               ( hps_fpga_reset_n ),                //                hps_0_h2f_reset.reset_n
		  .hps_0_f2h_cold_reset_req_reset_n      (~hps_cold_reset ),      //       hps_0_f2h_cold_reset_req.reset_n
		  .hps_0_f2h_debug_reset_req_reset_n     (~hps_debug_reset ),     //      hps_0_f2h_debug_reset_req.reset_n
		  .hps_0_f2h_stm_hw_events_stm_hwevents  (stm_hw_events ),  //        hps_0_f2h_stm_hw_events.stm_hwevents
		  .hps_0_f2h_warm_reset_req_reset_n      (~hps_warm_reset )      //       hps_0_f2h_warm_reset_req.reset_n
      // 
//		    .aescore_to_memory_bridge_external_interface_address     (addr_bus),     // aescore_to_memory_bridge_external_interface.address
//        .aescore_to_memory_bridge_external_interface_byte_enable (byte_en), //                                            .byte_enable
//        .aescore_to_memory_bridge_external_interface_read        (read_s),        //                                            .read
//        .aescore_to_memory_bridge_external_interface_write       (write_s),       //                                            .write
//        .aescore_to_memory_bridge_external_interface_write_data  (write_bus),  //                                            .write_data
//        .aescore_to_memory_bridge_external_interface_acknowledge (ackn_s), //                                            .acknowledge
//        .aescore_to_memory_bridge_external_interface_read_data   (read_bus),    //                                            .read_data
		//
		  //.pll_0_outclk1_clk                                       (pll_clk)      //                               pll_0_outclk1.clk
		
		//
//		  .hps_data_bridge_external_interface_address        (16'b0000000000000000),        //          hps_data_bridge_external_interface.address
//        .hps_data_bridge_external_interface_byte_enable    (16'b1111111111111111),    //                                            .byte_enable
//        .hps_data_bridge_external_interface_read           (1'b1),           //                                            .read
//        .hps_data_bridge_external_interface_write          (1'b0),          //                                            .write
//        .hps_data_bridge_external_interface_write_data     (),     //                                            .write_data
//        .hps_data_bridge_external_interface_acknowledge    (),    //                                            .acknowledge
//        .hps_data_bridge_external_interface_read_data      (data_in_aes_core),      //                                            .read_data
//
//        .hps_key_bridge_external_interface_address         (16'b0000000000000000),         //           hps_key_bridge_external_interface.address
//        .hps_key_bridge_external_interface_byte_enable     (16'b1111111111111111),     //                                            .byte_enable
//        .hps_key_bridge_external_interface_read            (1'b1),            //                                            .read
//        .hps_key_bridge_external_interface_write           (1'b0),           //                                            .write
//        .hps_key_bridge_external_interface_write_data      (),      //                                            .write_data
//        .hps_key_bridge_external_interface_acknowledge     (),     //                                            .acknowledge
//        .hps_key_bridge_external_interface_read_data       (key_aes_core),       //                                            .read_data
//        
//		  .fpga_data_bridge_external_interface_address       (16'b0000000000000000),       //         fpga_data_bridge_external_interface.address
//        .fpga_data_bridge_external_interface_byte_enable   (16'b1111111111111111),   //                                            .byte_enable
//        .fpga_data_bridge_external_interface_read          (1'b0),          //                                            .read
//        .fpga_data_bridge_external_interface_write         (1'b1),         //                                            .write
//        .fpga_data_bridge_external_interface_write_data    (data_out_aes_core),    //                                            .write_data
//        .fpga_data_bridge_external_interface_acknowledge   (),   //                                            .acknowledge
//        .fpga_data_bridge_external_interface_read_data     (),    //                                            .read_data
//        
//		  .control_bridge_external_interface_address         (16'b0000000000000000),         //           control_bridge_external_interface.address
//        .control_bridge_external_interface_byte_enable     (1'b1),     //                                            .byte_enable
//        .control_bridge_external_interface_read            (1'b1),            //                                            .read
//        .control_bridge_external_interface_write           (1'b0),           //                                            .write
//        .control_bridge_external_interface_write_data      (),      //                                            .write_data
//        .control_bridge_external_interface_acknowledge     (),     //                                            .acknowledge
//        .control_bridge_external_interface_read_data       (control),       //                                            .read_data
// 
//		  .done_bridge_external_interface_address            (16'b0000000000000000),            //              done_bridge_external_interface.address
//        .done_bridge_external_interface_byte_enable        (1'b1),        //                                            .byte_enable
//        .done_bridge_external_interface_read               (1'b0),               //                                            .read
//        .done_bridge_external_interface_write              (1'b1),              //                                            .write
//        .done_bridge_external_interface_write_data         (done),         //                                            .write_data
//        .done_bridge_external_interface_acknowledge        (),        //                                            .acknowledge
//        .done_bridge_external_interface_read_data          ()           //                                            .read_data	
//	
    );



//=======================================================
//	Turn On TV Decoder
assign	TD_RESET_N	=	1'b1;

assign	AUD_XCK	=	AUD_CTRL_CLK;
assign	AUD_ADCLRCK	=	AUD_DACLRCK;

AUDIO_DAC 	u02	(	//	Audio Side
					.oAUD_BCK(AUD_BCLK),
					.oAUD_DATA(AUD_DACDAT),
					.oAUD_LRCK(AUD_DACLRCK),
					//	Control Signals
					.iSrc_Select(2'b01),
			      .iCLK_18_4(AUD_CTRL_CLK),
					.iRST_N(KEY[0])	);

////	Audio CODEC and video decoder setting
//I2C_AV_Config 	u01	(	//	Host Side
//						.iCLK(CLOCK_50),
//						.iRST_N(KEY[0]),
//						//	I2C Side
//						.I2C_SCLK(FPGA_I2C_SCLK),
//						.I2C_SDAT(FPGA_I2C_SDAT)	);	

		
heart_beat  heart_TD_CLK27 (.CLK  (TD_CLK27), .CLK_FREQ (27_000_000), .CK_1HZ (LEDR[9]) ) ;
//=======================================================



	 // Debounce logic to clean out glitches within 1ms
debounce debounce_inst (
  .clk                                  (fpga_clk_50),
  .reset_n                              (hps_fpga_reset_n),  
  .data_in                              (KEY),
  .data_out                             (fpga_debounced_buttons)
);
  defparam debounce_inst.WIDTH = 4;
  defparam debounce_inst.POLARITY = "LOW";
  defparam debounce_inst.TIMEOUT = 50000;               // at 50Mhz this is a debounce time of 1ms
  defparam debounce_inst.TIMEOUT_WIDTH = 16;            // ceil(log2(TIMEOUT))
  
// Source/Probe megawizard instance
hps_reset hps_reset_inst (
  .source_clk (fpga_clk_50),
  .source     (hps_reset_req)
);

altera_edge_detector pulse_cold_reset (
  .clk       (fpga_clk_50),
  .rst_n     (hps_fpga_reset_n),
  .signal_in (hps_reset_req[0]),
  .pulse_out (hps_cold_reset)
);
  defparam pulse_cold_reset.PULSE_EXT = 6;
  defparam pulse_cold_reset.EDGE_TYPE = 1;
  defparam pulse_cold_reset.IGNORE_RST_WHILE_BUSY = 1;

altera_edge_detector pulse_warm_reset (
  .clk       (fpga_clk_50),
  .rst_n     (hps_fpga_reset_n),
  .signal_in (hps_reset_req[1]),
  .pulse_out (hps_warm_reset)
);
  defparam pulse_warm_reset.PULSE_EXT = 2;
  defparam pulse_warm_reset.EDGE_TYPE = 1;
  defparam pulse_warm_reset.IGNORE_RST_WHILE_BUSY = 1;
  
altera_edge_detector pulse_debug_reset (
  .clk       (fpga_clk_50),
  .rst_n     (hps_fpga_reset_n),
  .signal_in (hps_reset_req[2]),
  .pulse_out (hps_debug_reset)
);
  defparam pulse_debug_reset.PULSE_EXT = 32;
  defparam pulse_debug_reset.EDGE_TYPE = 1;
  defparam pulse_debug_reset.IGNORE_RST_WHILE_BUSY = 1;
  
reg [25:0] counter; 
reg  led_level;
always @(posedge fpga_clk_50 or negedge hps_fpga_reset_n)
begin
if(~hps_fpga_reset_n)
begin
                counter<=0;
                led_level<=0;
end

else if(counter==24999999)
        begin
                counter<=0;
                led_level<=~led_level;
        end
else
                counter<=counter+1'b1;
end

assign LEDR[0]=led_level;
endmodule

  