��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pi���.m~��*�+�V�[~�6B���ek�r�g]=O2������VH	k����γ�A�^�t	z�S6�S����,�8��`���7y�a$l_���n�b^���Lĩ��0�1���]-\>���1��_��g�Uw<`Y��h�~p1';�+�5pݏllDA����*����JRp{�+���Ä�ڻ��� &Kv^�͂�ӽ	��#5y����(�B��K�ݿ��#��-�H'�d��G�:9��>�' $=�xrW�LXR���bN��Đ���g����0��S`k�:����b�����$�g�&h��VS{vu�`?��P�!�(����o@O�����T�=)�P}]zq������w���[��PD�o�u��b(OO���dp��x�����;'���#M�]�|�P�����LSPC��l�޴����:����y�F�9����^�5(�3h��=��A�Cυ|ةD�➉���
+�g�|�'��&f���U�T����1X�2�7D��3�wV�Ƣ����`fj���]���(�v���$Q�6Ϸ�8����
�P��J��r6?wj�lYڿ�^�h���kKڎ솥�BS!����f|bu���w���[aT �#j�5'� .�W7U����=<y��; ���o���b�/iԛ�Y��a�M���(Cl$?Jt��p�-�v�Ͽl����X�@]��5
v�W]a��hmR)Ǥ�����fp�X�C�A�W�~�co���d�Թ@�joE�B ��]9tϕ؜�M�u=Bb*�	զ��g�E"ndW�O�Q9q��	���&[YĞ�O7�Ϣd&	��Z�����ɶ��FKg�$��_o;�θpN"��rP��!���oÜ*?E�3 �0"Xz~��$�'MT�θ�=�2�����1������E�(�^�EfK��[�|��Q������J�=���{����*��ǀ;�E�Ϗ{J���bL^dC���-8����`}AW��r酟�E�wt��/�_OT�R��9_�+�疱Vc!�������/������Lebbػ� ?�"��%?GA�'�,gq���>��|b%��{XjkA��0����Zg�$��Z�c�P[�y��͒��kc�Ry��>6e򛘡W�4}��逻z��3���zy�|x��=`3����������b�}(�M[�(��3XG��'��-���N^�ffqh��zo&�"�-h_�1n3c]�[}�M�9DO�}� �����?\��͊;��; (�(��al(~Y���}��6I�u�������w�oD�C�꧈�D�T(�d��#zة�MR�m=V�B3�2�^���.K\
�;�iɼ3**)G�6_��������3�B�(�����t��G��yx#T��R� �a�%�j�!8$�����m�3;�Ő+�R<_b�G��A0��Kl�nd��x�R�c�{�~
 s��M�������T���A۫��7�lx�y���o������ӣN�̢�ɹ����K�LHy��q(���&��E�Cn����v�wW��g��v����5ߐ�o;������_�"r��އX�n�0*���@(���	��H�[Oӯ�����$�c�xYǋ���{�Ĥ��!]�ؕ�(��'�rZ:Zm@>h=8�(T�=	�y��Ln6RN����[O�0얼�|��w�'/��\��ϝCw���5Y~����Mu[�Q590�;��z�|����ʸ�j����l���S��8o���R�[P��i�TS�,̡���.�� !��蜹����b���6�[n��ċ�@�it���̖h4��?���2������L��GaDRz�+��ߞ����xSN�|�<��
N�(
5@� �#i.�\��;�c�~~�)�M��z ��ft1;?bX�w�&�H���ߠ���T27���/��E�Ƃ��V�-���nõ��i���ܩ��rO����̑�mr��ZT��ޤ�vn���èɄ�3�C���>�Y��o�!��̸d��߿��c]D^��ю?�DYWg,lI~���n;�gYV�$�Өު��e0]�UC/g�[䴟�v
�b�hp��i��ޅr��*Cvߛ�-?
0-�q}�i�w9��|vp'0�#��FW��킪 pN7[y�S��h��Yg�L2��|L�")P9{��MQ�ߜ��8�v	3)UlOkY���oWt���z�C�Nޓ,�O1�=S�'�`nU+g�8�2���z��L:x���Ai6��Ӯ�rpxw��x]�[L�@�PR%H���N��B�e���:��X�X��]�\Og�%Ny��1E�� �Ufb�
�ƥ�'ƾE��~�w3E;���ً�8j���$����֊�sǂ9�I��R0_�㉕E��_��/�l�؁x2����(m񘌫�p�,KH([�$V������6ح5|DnmKwf���?e�a?U�/�K�j�Kh����7�U	�ר6E��a	�T$5 .?A+U���
]E6�����[zl�5���"1j:����D�>A��EV��k���J���#�Yk����mBL�}���5rΟ���E�+k���/���]����X�[O@�3%������*���x�'"�l�S]WpC7���?#�"Q9P���B��l���Z��hl|d+?G5�^�Ca�^`q�~a�-&�u�g_=͝�VT�p�������6}�jf[Q;0lpd��'�b�g�필QU����	���1��Cl��AuT���#����>d�1XEL�%��?K���Ⱥ�z�`?e�[�u��q(���Ă�$E�Bʰ1u���l���̺���A@r�d�\�k����-��2R&95��Ӧ2Zʆĝ�6^s �xO�Wu7^|�%qUt�����-wUw[P���OO����*�>2���_#UHޝD�J!��>f�Pz���/�^{�2���r{���6���3kʧY�����BǪ�U�$�෻^:E�N���?�\fz��Sh뵣����|t���( ���P`�
9�&��I`�ч�8�$OǸ7ͅ*@_ݮN�1żV���$�_+�Xƨk��D�!l�P�eD���,�%3���������J���@j<�~�Ӻ�&�H��j����·M4��d���J�ѝ����/��|N�8B=x��/����d� Hj� &{g6��Ҽi��aa����d�x�B'6�_�:�Ui4��O&|�8S�;��4��jt�;�<���~��>�������/<��g�*���+N���aW���x����0�r�"���0���b����b�����0c�mDrGtO/����O-��n}�
��{IU��k	����Rֆ�G�g�d֍�z�\VJUH��_Ս*M�)��d��:t!�ԇq�ا�yؾ���/���Q��f����	MSSR���!���i��P�@<lF��y'�0�`��;��nn ��&FFY���&����b!�ӵ��;�e�����`$��	H�n��v�d&T��p&�����j-n�+yk��'����J,)#�icԗO�����W���o֡k��G����]'8�Ū2#d=$k$"��v\����"s��9��ak�V#7c�M+�g���ۑ�m��0���7}^i�ځ��$i(��,�_I^ŷ������,SP^C;��@���O���9̙G�x���_��`z�7����,�"n
-j�F$RMY�c2���Tys *�H� �k0\��(�[�5A����e-y��j�2'&��L�΁ӣ#�L_P�(�������B7�ؒe��C�6^D*��/���,���(�m�02�����&�w�S��^ӽl���Ʈ��Ř8aK���LrKs��9�ժ�;x�N�4R&�g��L�)��~xzy�;VrO5!H�y�n�k �����?�Q���qhO���@��&�et4�����T �D�*��s�1�Y��0P,�^�8�z�3O�L�!UO&00����8�KF��vlK� ~N
ʵ���۳x��{�F����pVG�4����58�k�����]s���E]�� Ǔ@n�A�jja�T�FQ��=�7��r!D��XIg85N�B0���n�)����l*|lkJb9ת�3I�V��ۏ7*�\<������Έ�kw����'���O&����q����Ph��XtƙڃSu%Bq5�S�'k�h lOo�=��(Y*q��y�d�H���9]bA֏��HDב�S�_�J:�.����
Զ���5�+�=~q��[����Z+����nF�mc~��;��R���jW]�y�Ʀ?;�N�=���"D�jb(�k�F�Zs�w�j��X��TvCLY�}{�F�: j��E�&�ɛGD#<��	Tţ9~�@��������zA�/bڑ���߯��,ޮ��ܬeV�Կoq�jSs}�t�Nl�rR��\̗���%����Ȝ�����OJ�(^s)�ĳ��n��y��Q(=���g��ݳ��m�����p�����m@%3�KyC��x����6Jȓ�2���-�>$Ǹ*Gx��Fh�W�5��d�u�i��@�^p?��{�;�jb��$y��񮏊2�݌�]�B�R[���B���=�c_�p-�~9c�;���u����"q�� ������ag�����-�ɮUyx��?1`6
�|H�e�e��H��n_�pM/(p֖�eTR���(�`F��9xW\��X�01�ۏ��٪x��О �$�����ＡV��č�y�a_+K[��K��
�B��u��x3�R����oHt�������;��=]ہ[JzVC�ٚd9��JQlo<�8��ep�{%a�e_���V�9I�������3�P�z��{"Ge�xZ�7�EЎ�a3O�ʶZU|��}���`q�����|�x�r*��/*&m�ڢ�aA�˦����l��]���WU?f�����ZJ�[9�1���"�]Rޱ��R�R��-�d%@�y����C��|9{�8��ʞW����À�x��®D��_�nL�_�T����.��<B�Z��r�J��ݖ�t�V�M.��f���v�Q�wLMNZ�Y��H����"��me=��PJB�N��tc��]��M��¼W�n25���vI�����?����e��N��g_�F�hU�{��Y�L�0��sv��Baqi��9�b���0?eA��_]��EB�U�K��XV�5Ī��֏�ԥք!0��
��Փ�M�yp�%_��X�SEE�7�ӽ�oU<A#���~�|�
�&�#ծ?��S�5i\NثZ$6��˗�[�"f��{�!ޓ6� V#�+/?;1��p_(��ݹ2���8!lGv�l:m n��;<n� ����"�&����̳ƃ	Ml,&�GA������,�U7���&�*�gz8��Z��wB�aކ�SS�MJ����ǉ�-�d��K�o�7�B��/��&Y�l_a?���P~&%T\t�QRy���It��6]O��!��D�3�3��sn��I	�)�*_�^Ps���T�� %��B˫�r�{�b����ab�W����l.kJ�9�@H��g�ܾ��x| jV������Z7��=�e�)����mΐJV��	3�sC��
.d��pz��I�[,�D>�����sD-Gҽ�u�l`H��C+�<��l9͊L;�Ϩ\J�m6vsoU:��������F�YnhJ�䪉����A���h��6	Zds��\M��ޗy|��kM�L�U�I�z*
J��+
y����Ф-wi`�P0��04F[������k�;������^���,�9_����8gP�s���J�{�	�85ͳ�=��/����غ{Z 2vT����G,��f�(��}eAU�YaZmf��<"������,���)e	��Օ4ǝ���A{-��*���pr`֒Ix��w��Q���4�Am+s�.��ϑ�TԔ�����uS�|gx7#�baZz���g�N�@�C(��E��B�5v�(V3�m�4��=^�D6M�cD��[豚E����S���0����.��Lכ���D2r��ڏ-C�^Qeg4$���J��=� my_��ዓ�R�s,����÷��ح�s�+�� ���C��3�7k�2����_��T�k�HPh���r�Vևyt�'���b�oK� �Sз|&�7�ዕ�I�U������k0^���he����:eط6F����'��t3(9h��cC��|����7���u��<�S%~	Ybx�a	�,����6���$����n?�2�\A�g��令�)�Y_��[Z�Xn�΍}m���)+�I�~�x�w��F�m�pm�7��{BW�%�RJ�R��Xb~S3��L�La6�&����+Vu���D|��-���X����Ę�~����otW"E�QA)/K��N�K@UeuL��"�i�N�/z�M�٧$���Xe� �y})��T�/��}=�boCN^`դ���Ň('w���Z�{Ri���|��@�8�e�����+x+K��t���÷���ɺ<��|SA�ڢ*��K��Y�r���ʹ�c6R~���&����"B1 �_JvWt��6B���A�M�ʮ)U{w��"�+t�q��3��,o�&�Wgr����d�u@E7H1?"\�V�ڶ~K�g��Z3�E+7�p���l��hӢ�0�Y/<%�  5�vWD]c'R���F��Zv�K�t�CӋ�4p�SN�&�I���Y�C*��������{�7����+�Y�_z�n˼�b�a��xw?��aQa�S�����R��� eak@Ǆp�� {�\Uy�� rw�LH���_"�-U�9�Au���p𷤙�[�����I�|�=|���Q���fr*�?��nl�r��5V�8��G&n��:�e���OРЮ����9��3�e�@���G�<�ڥ׉�;Oˏ�e��G�ۤt� Xv�޺ZY���w/�hZ�w�0����c1�_$
!9Y[��}=�X sdڼF��m��K�x�*m�N�A�*��%|�:sw�AT�̂�˫q�Q%s^J�Ԉ�p�xW9�@�� �{+g�ɿ4�=�O��%z���&�eT�Qo�V���%砒�.9�\MS"S�=�\n I�3�ڜ�)'��b��Ew���C��m�5��KY�yr#��g�>��cz�3��[���f""�C����.$��9֊������Z���c:�Ob�zg��.0�Ց�Ĺ�>1�����\c$�5�ʥM~�d�jN>^��B0p�`�돣:��yt���֍���W�I.d�����ʦ�� c��@s9���Oq�~�u0���$=�m�9���du_A�ѧQ3��~Ur�xB�!�����3�ׯ�5��&���{��&L���D���F����@�Y���c�/Q�#2j}CR�����E�k�Tv�UG�бh[	��w!�����ԫ*�l5}�F�I�J��*h9ͅ�2�R�2�e�4ڎT�M7�2�$�T�pg��1�l�� ̆h���S�@��59L��i��v!�������ض�Ag�5Km}\�qkC��#�}�r+��:x(��1rQh��.	qI���`��kVfR��i��AtN�ż�b�(�V���_���Gw�9t���Z��Y�Ʊ�|$��=֙����7���\y��kJ�K�����z��,o��n�3^��L�\�2�̴U� Kb?!i}��䌳V�V�B�.�}�3�ņ"L��I}-��뫈���
�J� ���`��C@�H�Qp�^�̀eE���B�c
����O�4�b�z_ljV��N_�Q���J(���3kw�ހ�'M�Q>j�<tg�R+"^���=8�ؗ:>퍡}�,=A����)�%z, J��x�P���Rp.��֑`�^�/a�Z�^MM��R׈ud� p�U��1�_�%v�/��#�H�n2�C�_�&I��6!"��P����!p��·=��Q@���rA�gh��ߩ��)S���m�i�'�0�=<d��/�$1�Ԙx�L�Wx8�3��W�lxh��c$�.]�ۡ����U�@����M���ڿ�#�7HP���w"1��	Qj�"��-B�f��Ҹ�y>��Di}�$�LuAN����U�<��G�R�������;V!e�i/��}���	���15d�:I���.�Z�U~��Xj����iA[���5�F=�W�>Xd��EeҲYP�N�i��}�TkW���ӭ��L��{2��-vj���4aZ���s���0d}S�����m����`���.�k�Ud�&��^��YD�w�Xb���X���'���Ζt1����@yly��GS�\��R#$�[���,[�jV+�Ү��t�;S�Ri@V��1+s,�&�����[@ًmk�JW�ۧ$��f��'��Q��%J���� �n�6����̈�]3\6���!�����7����_�^-�^y�A�h�3�P���s�%0{ދ�� LD`�%>,�d��K�$}mw��դAdJL��J�j���E��xMpY�VY>f���'�&ǟ|`�\��^:?!�"�0{]� %�U70��>�v���3L�|�r�g��G??��@`�VT�g/���h�v���^e�W. �Ѡ閞 v��m�0�X�-�P��M�@����,��� `��O�<����:�F��h}_�JO���*#�C��JH�g�.�t��mݏp%eFm*)z0���I|%�_�����Ƒ��l��_UVm����ř�fmp��/Y��b|U�r�c�SmI�X4if����\h��`~�'�e>LQ��޳��dwܮ5E	ص��H:IO���;�$�y�����m=�����h�|E��"]��g�Ņ�N���-Ś��e�\�\��6d,�t����Y�8 ;;~�������md�]n�Z��bOY�5�
�æg�4yhRX�9�G��ASu���EN��|�����,7�f��V����1k#;ҿ�aC�*	(�(C�+�ܝa��N������)'1�MT�SZ�EYݦ5$K]2���C�["ʗ'Mm�����g-�l�0#"3�\�2#��t� ��4Ƨ76�����,"'��`�{��������ˆ/��zR�����ve�B����6z1뻽��1k�*8L�b�'�Qkf�z=r�_"����>��d�����p�����B-s�b=?�ߛ?�Z�nɌ���� ��� �m̀'C ,ȝ��&�Ϙ��*x�Ȥ)W���n�l�$����D�Q�U�?�A�V��]2���o3x��}���L�o�S��ћ�p
K�m�d2�2��S���H��X����[�%����w߾C׌H���R�<z�3~�w����S�q���0�6��З�����ޞc"ō
�{��^�-Lm��M���p��'���Cm��U����6<��*��j\��ĭ���H]���j�0��(�����������X*��������˴�U����PF��^����2l���+g?�k�1]4F��(�9��X!�U�ې��L�u��}dr����q�ꖣ���Ia�{;�O��� Pg�#��v���\���`����m�Qx�E0�I^a���Ə�Ӧ���~�v���,���Ĝ�Yh4�̩� ?����`���VQ�W�:�0�;ZI��om�#&i�����<5d1��Z���6�9��(6;��;A�_�#l���A�Q���?ԛ���T�B�Q��q0z���eMt�ֵ����/�.�e��$O�[�kn�r���qjt4Ō�:�;<�5��j�E��<���)��e$mVbV/��[oGt�ζ̆z�����׾35��V^H�A�`� �g��L�ϟ���Ȟ�0FC���*�2Q6q4a?���%�A����Y����U����8nP���ϑ�r��Q2���|�q4�� ^�eh��c�h��o�W�;4�F���~���m��W;�|�w�7��*}�VN�������v"����& p d�`��5t9���pͤT@������8Q�m9���Ȋ{�fEn���w<i��&.�t��z����UxOh�<V�N_*I�}���Й�9H�r�<)Y��L�wn�h��i�tw$�Mz;c���� ���SV(ƈ,�NRB��G�V<�-���9��I�5��?ȟ��ʻ�^G,�J e��'��v�G��FKb&�n�1�?�t��i��=�ߞ��F"e���2�f*"w������j��c��7Ie����,q�p��([��0{��6�e�H�Q��mo��Ș9MU�"�Ip��ۍ<g�˝aj=5���r�0�Lġf��Vg��r�\s�鬽�j����6/8_�:Տ,��'��K���7�vƝ���k���Ʌ��N������2��m�w��I$m_Y�8�-QQ�y�9�:˻Rz���̽��k\ڌ�����Mk�c�'")k�lt"p��z�8�|H��G�j+��M��T�ϗ�Ho0��1�Aɓ��#��&RS@&�%��^k���d����(tY�Ƹ�Ը�~Yr�����JL����g���m�Ո��esz�4�*G��C�WWd���,c����+ܧ7����['��k6�hʴjP�L�!$=�*��MZ�-��3d֔�2���aCx��m:�!D+�%�R`�b�K�p0���r���ѷ(býz��y��=	�߆j���jUu���^���<d+!�n�jaB��uԸ�ҭ?G�����j���[���G=<�&��]K��I,!Q�xP��� ��1`�>]�O=��MC��q>8���?`�N�2�a]��Ǎf�3F%�w�*	�:o?+��Yx�gL��w�8AP?�]s��7��Mkn��+��R"e��O��h�:���k�5_a�C\�+�b�7z���n�?��_����Dd���A`]�r��1�m���**N+]�Y��/��K���ټ�p�+<����ω%%�����I��(�:*Y �zy*�4Bn��S��ђ\W���m�ɷ)����Pv5Sl�G)���@ ��t)u�+�_[��#I�f-+D�;'�Hxb�'��bT�O���Ξ��p���&����Y��'�%�q&S25�$��t�*�jч��!L�̉��B?�
A��� �PW��E3�ڛ���T�M³޼0Fdl�v������X@ ��G�$��W����������Lô�9�4��j�(�Z\!�X\����Wruo!����]I'H����d��=b"QJ�g�II� gs��N�g�(��X�JwT�@��(cto���`,��K��bc�LBxH|�3Kf뉉o�U��z_�=��X��Ii8���p	[���m+ٻ�,��g+�C��N&�*��u^��n�d+�����(�V��u8���&DyxK!�S����tEwԡ=��W?&�f��$U�'�+Ao/���ٽ9�2����0�\�Xl�SS���ֻ�^n>o8`�J�*s�Wˡʿ�5`�rD�F	5[���P��GA�S�Y](��o~~-��=ʝ�p��~�Re�B��
�Հp
�6��gX�_DH�gq�����Ԍ�pW���)R�XY�G·[�J�I0w�Ȋ�s��.;-Y�ݮ����vU6����/l���ϝ���ع���߀��	���Z�m�C7�^�F�N�z=!��#��e6p����unt�Q�eM�e�v�I�����YP$9 ٕ�)��A�?yA$o]D\_�;s��fP#�UQ̪u��j�5F����Λ�
1�R��ō[! $�5ԕ�O�+�=s�cO�LcI6���],җQ�z}���&-���|��zL1���\�N��ʉ'�Gb����E������G��Uvl�B;�P�O-��lo*�c�����8 �VZ�Ȃ2+���.�'�����m"4����Kv�c�~���Ay�W*�C����Hj�1C\�u�jd�:��k��G�44��i��Ct&�#\g�Z��)Pqtf�oy�?fEȢ��٣'?B�*־�s���AFc�C}�Y�W�Ȃ�A*�9���a𚾞ȋ1��"8E?��ˬ�͆S��*iCϺ� a�2�H-�@eg�=��M1=|�ۭ$K����7�Y�I]�/�5X����?�4�sN���y����`��p�:���Y�2��_����@,����>r�8���:I��?��dz$ti�L�E=�"ib�a�`�<Z�T3��?u�C�FV0�R���^x(��3��h�Cy� 8���°�z^N��C����f�&�sَ^�z�v�y�)��e�� �<9�����1=��������6��j���/�F'��X�`x��:_c�Օ�u���!�d�%D�v���������xL ���=:�����]��yt� l�t��<4��z<��Z�;#0Δ�.��߃xh09��y��V�kӏx��	hI�]E;N4�˙�'}$E�g �X�?oq���͉��0��	���d�/����.<}tNE����m�)'����z��,�/�$�
UT�	�N��\7�xQ���a^4#3 6|�6|�;��	 SyZr�L��V9�* Y;9��i� {� ���)�&pW�n#.ɂ�㻝�r�Wq�+�8OB݈���o��4)�:I�n�K������U��[[�>��R��MBjwй���h�H�l��O�h<Ŧ�{}��V_�Y]�(Jn�R��qJeykl(�c@����c�ƶ�~ɏT`���g�Ijy]K��E��&O���ad�5J���A	��_%%��y&qkӊ<���ɐ��_/o�uݴ�!H;\����@���g^;��6}mNsX7��V��Ԙ5�K����i}�r���:3���Qmi���S�]���)[2S�pL!��ڜ�v�l���8�C'ao�"(������F�@����0=nU�g��
6������#"��x�f�he}})�Kݐ��Y%� ��X�ٍa��cYc�S~���y�������Y�эV>ҩ	My�����}9ٖ�('��B�f��=�2G���g��u9'B��f���5��@��_�:�����2�v���@^�1=�{̉.q�]/e�#o�8�plu�����F��M���w��!�Rd�%Y��BGt�7����u�������f͓P�J�fF�G��
3�--"~��L���땟�6��P^�f�
����G�k���ޢN&���D&�^s`Z7�p,�i"�"��<*�J�տf�� HU��pޒE��"u��=��H�R�nH �'�)��=��+���[�^�mYX��c(�/�X����$Sf���vQƖ.$=ˇnPh9�$�eRe�䢇0ٜ�$0i+��s�@]?�(ph�F��J+I�_��)[I�T��P�˻��5���`�U��՝������⼋᳟b���{��@�N����<f�J���P�1	G|
�Pd��D�q�1�`ʍ5�mNh�A��>�G$��l�ccl�Zf�3������ �Z�tE�D�)X$Kfd�x�^տ=��g��v+�_��E;��>���v�4���*:}�aⵆ^/EP�>�̡P��Me����̤$M�+�bH�ڢ���5�)ҳ䶨$�&���D��N�X����zn���H�E��%��	 J���}
r6�ٞ�eG��B8I}詢h.�m��/�F��Nvx�*�.�Krd��6g�>2��fE �k��w�x���`�IYf���
mϪ4��5������̧^ŀ7\�	+wr�&�N�tA\8��$��S���4�P'��V��ge�y�?Ne�k.Vgz4��Ba��a��i������;�P����Ubw2���Ӈ��a��4��6fo����k^��n��?T:��[U<Ĕ!a�^�{i�D��{�%Z:�"�9�(���GІ����>���,-�z:P�k�H�����Ƃ	8Xs�����o!�kH:�\�c{ v��k6����Fg|:D�I�$\���N���١��jQO��HZ�K��ߺx.B[�n+ZmbLD!b�y��>����EL5}����p�ݬ;���x�~�/��	���,ά�?8bI��߃��f���in�G���� o�A�aas>���Jz8����*�v' ���kЙݲ��-~}�G��[�^P�"���L�5�$z��M�7�([�D�[U��>��%�?�}P�i��4�~��Z"�������ܮCb�)�^��Pm���əB,)�[�;���+g�1��]cq�,�Ik�_Bν�B�������n��k��ﵵJ��!������u�u陕�b�dZz�B9'-8y,�У���_m��N9�4�\=%Q2����	Y���5Punj�H$��p����H�W���A�E Xr���\��F�~��JZPM0���|ର��U����h����������L�����[���4��2q��A��a�W�j�^�罿}�eufhT��|Is|���2�ՂCfWqMǠ�儍�DN�s憎^ԌA��c'�y�+͵��������~L�(XDJ4%&�xg���A2�|�w�9;+�����M[���c�ċً��!f�l]�7��]��ڙ���a�)�pҙtW|��	i/"6�(��al.4��/��z����t��a?@"9lە@��>�ij���m7��\�C�z��¶߯��LS(�d�w����(�|�x�6�c���Xc4������a�3ͤ����Z��??%���u��#>�(��*t����s��G�GQ˪��2>ͣ��~h��f*|�����e��`˨<6��
��S���lF�V%�W�m�K�eh�aֺ���z��5���I��;)��W��y���/��Kt���M�mA'b�O� ��,�Ez4Z���3¤)��y����rD�Gl[I�-߀.��rY����6k�G����Y�~^N���G!��B�:at����X�����B���{l 9�M ef���O b��t9��QGF!���Γ�xФ'=�p��4ڥ�b%~�<��~1s�7 Jh�����;��NczOS�l �.2�3;&�$�