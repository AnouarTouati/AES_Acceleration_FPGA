��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղo�(��3mM�,F$g����]P<��=��bF��a<�Ғ��E�|+7���7��UxHm}��4)a��\�CO@([��\�|@����Q���߆[���C����]=}�J�ٔ���E�*���9��2Vg�b���Սk`]m=����7!2h���]n�%~:��(L�I~ta��'yKh�4� ���?�\ِ1�G'I��6��m*W­�.(�A���Ԧ�?@ RS�GRF�ީ��&�������b,�I����~��gD6�V��`�S$WS{��k	>
p(�Oh�P��|���94���������x{�V��Y��r��$�Ӡ��`B3/V薇ޥ���@iOI,�$���{I����X���/\�n���{��Y���Fȫ�d����kc�졁��ߑ$�=�8=��ƞ���6�7|M�"��zk@oHo�$A|�U܂�E��L�Cs�ȝ����:J�Y�d��5̄�����u�-�?�;����:� �p{D`��M�7N"���A\P�=�Э�Nڝk���*D:�9�P�H)nS�͐n���q�!�?*	5mk������(㞔���;I������;|ٴ����D F�ш�˞� ���Huߔ�5Q���&m��ա$�A�.�f�]3p���ng���:�K�57mD��!��m�X��p���m�����(�w�h�@6p� �����"s����Wu�<�r�@D�u�b���b7��uT�I�+�~�v��Y	�H������#+ŵ�&7��5a}�v��Lz���L�?�'���72Um�є�����پ�a1�L�..��~a�2d�g 6#H�	<��xʯ��w������DQ8C]y��A��5�0�-������Ҟ���4<S�r��l�i�-��>����1��Z&�xj��+o᭪W��4y�B1�8V��ʻ��)Gw���h�E��9�s����C���5��rg�$�i���݅aM�`�XG��D�+����[��lZt���c:΀��
�pӂ@���q՘�*��J����ۂjVf���X������}�@o��fy�l`7��_��u�$�UL]Ln�nX>~@|��!���y�#ؚ{膳ꍆ�w�<�����6+R2���~�ł��(G���a��\����l��~�	S ��A����Mg�
z� �Nᚉ��΋&����-6E'���i#��w�ȭI�T��:1s$�DX�P����N�Kˎڔ[F���f���8_�G>�'Ie&���j�S�������;W���= �˹�%�Y� 8�1_6Fw�]e�o��ޯ�z�o\�d�ap��k�ܐ� \�J��)���,��<,À1����!Hu�fw�A�-�C��I�0�E���$�� �{��(}�y-����=~� �U���铮�ٜ���P���`�	߹�!��
U���Ul.J��߿�\��3i�!<���ۈQ�Ɉ��V�/�h��2�72�E����Rƻ`��7O�����t��?NpƘ�~�\��m�1|9��k�� ��HAz�'���[〔��$_�Cr�S��!�tD�L�\a$��\l,��H���������� #��9Gsq���d�H����I �<�[���1�J7_4p��*2�C��r�>�Ớ�@�|--�{b�5���˞c��fW[���+jsݢ�g5��������ǵ;�r�Y�	�	�0�G @F����	���R1��B�,@��-a�I@�>#h(o��=�,z0ЕmQ�~XS��/�\>�/��R{�e��T.�����aݙ��?�MՀ��?�0G5zk8��+��9�B�<��x�W}�+���� ���6;]5�i3��ʤ+D��kc�q/L5�9�a85F�G������y��@I#Y4.c�D%�D��+3����8�'X��lTέ����ԍա�f��DJx�Ͳ��Y�f:X/�쨊��W�^�Ϋ;G/�ɔ5���8/:'��c�ZT��Zu����Qk�z����)��P"�ᇿ5�P
������Dǅ��IC��;P@�E��kr��2hv@[L�%�N��� ?�ݷ����u��b��yfz�@���$��@�C؞�Ľu鑪z�M�pe�ò��$���N=�ρ��f���()�^Ywo}��������z�=rJ�{p������&����I&`xu*��M�h'�^�e$"�zS{U�9}6v�D$ax��P���q�����(̯}�ց"G�޺�ٖ

N�V
�O	]Q	D�r"`��d:��p�����{�p�K35N]��9dy-i��3,OU5����&!��8�j:s��/�^q�F�@�s�,�m��]�1 ���A�'j6��o/�o���.w�FS;�
�X��3Lәp��#�@<l���{ϔ-�����R�fv$H@-s��%���<�Nu�K{xc������n���N�؂�x X<5��}��M�GvrWEq��P1�z��Իq+�S0�\���㬷����Y���'�3�����
%� j�9���_�� ���N��|�?s���4�?2�>*K���b��ށ(���f�r�Y�;�,�'��	�����5��U�l����{�D.Gev5$�s�Kz�u ��)�t	�iKc����͘��fbDJ��:����<v�+��*�?�s$羦�6���#�"�I	�[!P�V{6���&��ܰ�\Mb���<!��z
 zCo�P_Rդ�3x���ߛ��|��X�;�z{���A	UUhǘ<��s���Y��f�SR��"x��[}\1��잲��dK�3ґ���*���<�vQ!�������^c=�Mw;9G����Jf�z5�D��r����;�P�H�g�4�\p��d���& u��L�)�ٶ3�H�Ѕ���/B�&a��w?��������;��ڪB�M���SF�=���5;�۪�n[��W���H��]�c����G�ʻ�>���0�py�R.ALf:�zĻƊ�eȏ�&�Ͽ��T��*���c+��eŗ��ƿ���G���4��.���g1��WK�\���AwK��<�s\�_Q�l%a�]�Õ��(ܩ/I�x7��Þt�_��?~�a�7�;ƺ(��ѿ��,��g�ő���mP���4���G/�58��@f,C6j3""�*Y���:��hq���]�9�����]�����=��Q��?��qӤ�&�*Q��{�D��a᷄���z�o��Eg&8u�|t�=����:�H�ބ1�h@����DI��,�N�>1��Ɍ��Ō���p،���* i�a�6������-���e#��7����o���
�c���;ٟ i3܌���%~���C45<��c��4����ͫR�i�Q�;�'�/� R�\�D�l?K�F��^8����T٬"�����9����W*JTyM�#G�YUk�2�jܗ�eh_�n�e� %���"j����#�#z\��bb��(�yJ2p#i��
9 Dn#9]�К��y���,��%/��=�'�WC�jG���<M�$���@���LDd��i����O@d�u
��|�� Ҧ�� ���]ٿ�BbAA�m���,�5G�|iJP�=â�4��4j����0!ж��(D�꤇Ph�}�{ŏ5�8@��=�"�[���Th��V@.�h��۰�i�0�,��rm�͝�&ؖ�Wp��}?h�ia�9���)	A�@�k��hڷ0ѓ%��
����q2�c�>Ec���eakɀr�����qy���*�L`�Vg�/�Ko}������;Ir��p%��	�.�sq?Ӱ�H��J�.u��/�E2��-���2t����9�@H�|��SmGCC '�୽Qyb��E�����}�\=$]�}�kE�811����؊��IbK�S�F	T�� Vyn{f|+���yP�HȂ2��Q���L8`��6�Uh�ew��ǬT��K����I=�P�*e7[�� �$��U�QIR��i����Y�s����IkWF�[JM;�;p���R`Xe� ���#X�w��eD�?����7Z��&�n�zJU��S�4�?��T�5� ���d��S\ ���ⅈ�_��8�n���z83G41���"9DJߥJ�r��ٿ�����0���Qk�2�[�ѶM'��`��|����&��a���a��Jܥ/v��밌q� �]Ȳ	�r�́�Bω�A��/����iYd�O��g���R��4���)U�9ĸ��!�S�*���5�V<\S8�i��\���`�/�X2����>�Ft�hU����/���B�z~�'�XW�����j�w�^�)0)Rc��읇ى/��͆|7�G��&�}CeeC���Sq��
�4���BNf�����vZ���\����C�R�vTL@C����L�F�]h�yà�/���Ńn��o�}�t!���W�`��U�	��w��6�eSKZ��чGo��.?ߞ�	]\�������Ju�V����*����C�nR���iz�\��v��:Ы���Pf�{����<T�<	�����B9F �x�� ����9���CQ��OjJ��F�׀�ej\h��/� �\��XY�Yꐟ>^D�R���Cq=<�z�Dt���/Լ~SC���+�6�賬7�Pz��F�u�-���Ӹ�fm6�/������vJI�צ����2W�r�#-D������tdX��`��׆Iw��^>y�Tl��I���J�[� g��Տ;�"�1���`Z�����T�OY�kL sfp����wU��d<T �*o�����D�&��M�է}�ba�`��B��6!;��-p�?���K�_�*��f@�������c�@���u'
�h�ZU�<Œ�
VP��d���3�@C֭
Ku ��%�������(~�\�z���pO���.Pnqm�@g\<�Ȍ�5I�y�B�� �"�bi��+�֯ݜ���/�#!�d��<[s�H��g��n��q�� ��&)����H�-}]��	�f�vk7��Ƹ������)�����V��D !o�ԩ��
,N�E��!��0�{ c�ҭ_.�3��<���K� �[T?�4d4j��Igǩ��p����u�:�gD��)N� �j��{�C j�0~��r"N��uѭ�%&�K]�!�Z�"�x��&Sm�8�H]~��
�d~��6����kd�ߑ9�vP�Ў�nȚ'*���Ŗ��q�R��f�
X���������]"���lb���Cjw�#�58ZsL@�:��^�J�ȴќʀ�U/5(d�К �\�>�^*/�zIwo��$�&_��޻c;h`������2|��d�qL ���n����<n���vSM2��h1��@º��۞tJ��HGPzlv�ut���̫Ճ�2Er�;.��":���ק�%�C����m�4�Ϟa=�l��Ҋ��-ȕ�v�p;7�;�-�y�3�4�ꤍk}:���&y����5<E9<��^�,_d���K����Z�� x��K�MY"Ƨ�9�'��)s�>#�h�^UJO�V��h!/F���J!]��%>T���ܯ�Q�L��7ჴ��|������
����[����j����L�hz����[!�{ZG(r���Jp���e-�B���&����,��ː}��?FȐj�3�`�nan�ix�3���u0�ZYM���R�fgO�N�D�<����B��Me���ӌ��K#�K���1$�fN3���1���{QRE�s!)k1b���dk�Clq#K`���8D3��s>"�\���2+=�2���@߽:�k�PKhU��zȍ[��绮�Ɔ�e��Ui	���\KJe���%-Q��>�ɾ�u��,��UM�W��0*�	�hB�ߘ�r��O?&�~I6x1��<�-��$g����L<�w���M����i���+�������P���t�¸Z�9Ɛ@{?xn�=���CmvT�C�s��a�������S�n��o��ߔ���ќ�g�-uL��o�jyUD��w��?�m�3�'-��TJ��!����K��K��S�(�|��QM�(�6�E��#R;V�g�{Ej�T�ɗy���x>V!�̯�Xg�˜8ɞ��|Ѷt|~j$�S�i�D�=5��p�E7ɉN��n�k���M<KE��<���^>AZ���Va��C���( ��؄�4�a�GS-�u{�O�X��
�k�V�g^�ro���=b��*ǳpA�"1���G"f2q�T�\:��%��e��]���qӡ f��
�a��j�q�x��Y�тu��АW�!��>!⥌U�g�r�$��>�%��\*Z�����Cqt��\���A�Bi��f_�:�3��EE��ׇ�����3ͽ��K�J���%��H�#!l�#�3����q�����&��0�mk.<PsΑoCF�T��k�+屹�_Ѡ�a�@a?����pv�}3��U�2A�������b�A�/����0X����UP����#�z*y'O�y��u�߄@�@��-��E P%�����e�)�E�]zΑљ�|ڑ�8jdFG�+7f��%�r��"���I���Lc�?:�3L�1���������$�
7{l�}�mh������20�w���Z�Hx���$�no4-����dм��m!��;��l��C���3ned< 9#'�`�4����]r
�I!r���I%"���S�!����2cqՑ��+����=�i�����)64;o8тf����Ф�z�֫��v�^�����K�"Q�ߴ�X�`ȵ�4�\�;d�*��,���4QO���ۋS���Jz�G�K�aK��,��y�M�O�>�o��o�O��;���X��y�k�_ĺ)��&�@��+��*������lF&a���4]����94@4�*��&z�#[�P&*%�^��ՊY� "�|��Q&��F_z�%(Y���E[�L﹂?+��7у\|��nF ��"S:n8���gAP�����n}��o2sع����mN0O�o���
Uߘ)ɡr<���m��|P��G���F�n�΍�;�i�5��d��Xj	���5:"��h�4н'*���/k�����@.sqzy�[�$�o�F�ĕ�	��
Õ��1�������"%�\�&���.��p�ϋ���\��D��60�*�Zӣ��`_�[�[�p�	�+��IU���I��	����zk����H/8�p��C�XL���w����G�����i�𧗏
�<" |"�Y�=�M���,�
��x�C��Z*T�AC&uGY�#�K@����ƴ��F���,��MP��BE���Iθ�w~L���/�� 	��H%��[ٚQ JA�l?.��i���;���~j�[&�W�6LLĄ�B@�WY�����U��D�[�?��28�Tav=3x;�)&9D`u'�<1��~�@��^$V�&O�F�M0>����k�ɛ�����Q�h��O��^��(��"�8����K���@U���>���b��)�t��W&�Z�x�Y�5u�$M��Jh6-!?agc�Y���&|��Yp�,���2Tw����Q0��S������@I��4����M�;m�c�s���+��@y� ���JJG���غ|A�S�$!�����"�����kjB@���M�_��=�J.H	L��9a��P��

���~���V������_h��jp6^�&f#Ns��m	{�C~�;�"
�ڿ�~E���� 碬��|�M��l�&?�,Mz?�dPoO����gt�;}��չ.h�\%�U��18����׭x sK��fa�|�CQ�;0����C_<�]%'mc��Z�_e�5[$�{��c����R:��nӊi��x/�	�,��Ő�ڇ��t�%����s(:	ු����<vz��+,�@���8���N��ׂ��@��:WY��� e�I�y�Ս�	�eYf�t���+߸�m�|4Hn��y�Z]N�d�%��p@b1��/�TXڍ8�faL��q_L��A���K�b���h`ٞD�3�bG�ӿp
��Œڪ��f�B[��(�GR��~#�
�~��gZTS����-��VM���';����.4}��S�B���+�3�wb{��Io�����g��o�2��`���;�Jsނ���U��Z�vQ�r�h�u�/�eU	��J�Q	������U�hQF�еU� O��e� ��F��ٻs��BQ��4�E������Ӛ�v�&�v8R��r�6I�T~���ehf@q�~S,w��,Ϣ4�ᵗ�ŚA�j56�Դ�$4]s)E���{�� `���!��0ֽ������F-�{Z�*0�>�$�,s��L�G�.J����lĦ���M�W�3�Yrt���ԞR��jӢ��ʅt�!Cu�BK����6&ڏt���R}��hJķ�������
(�Y\��H��@��@���\�.Kk�arX�e=*v�hJ��T����0�5�o���0�� �B��8�r,����z��&�C<h�������܄�NQ�R�Q2j�4o��w���Ōy��%�w����&�`ʘj���	�٘y�T���K�i)����lV3,��>y5K�dTs�H�<��T��\A�u%�ת��ć�O���?�RC�����Nϸ '�N����V`�}R�l:�35;���v,e��l�ex�`�Lv�r�1v��w@
�m���BB�pJ���������`��'=wVM�&	p�p���m�lR|�w��]�����^ݬ���۹f����T���Ӊ��6=�r�X���l�h�	4W��U�P)�����3���M�2��(<^=�o�a+7׶�����7�f�;��L�B�T���'	n�n�i�����,�����j���
j�J�沺�d��9s� ��n���L���ϣ|�w����%ɎK����Vōܾ<���Ж�4��K� ��'Vx�3	(�9���kK������_|�4^�����Cg������#���d�Š�Z�,/�c*ѽ�d�g߸�w܀j���)���U -��0:B19r�XU�n�#O%����Ng��\�"�����ӽl�FG5����z�(���/qV�%Wۀׇ�!w�94�Rg�r��O�A4�c^�X��吷�@^��T6U-lԛ��]EHnֱ�fl	k����:���lk�/y���	�b[�?�6�o�uJ1��5��Gi"�{��5�"�F�^s����y����v�uk�(��r�����@��i�U����=u4�9�ъ���ђ*�bP����՛�?�#���	�Yt�%[���|���Y�!�7 ���;H�q�Z�����]���/)`[��J�h��4�a��\ݦ�a@bu:�� ������i�j�®9Z�oC���$@律gm�����zl�M�u����7��O�S^�y��X�%230�N��#~�R���XbQ�W4�q�v!6Iz'2u�;=
�|Ţ���'����:Ѱ�غf+�����Ô�a��cn�5�7��Pɛ������)��$p*���|�
���\�4Ք���Nk9���M�7�����p��\�j�l�'Q�����9
�{A��L�%I�~����㺁--V���B�w�a���9�<�N��� ����o�0OB�hW��T�E߆_�*�����[�n�%���G����T�6�"�������GQi䀆��ݯºU�(��4����w��48pY�;�N�8��9��o@_����qV66Gb.u�ބ08'�5l�L7�����4�lp�/LSQUG�E�MP��kx�z{��j@ XdX�v�t�O3iY����ʹ�|��5:🠴b�����d,ß
��Q^�#/�cK�`\���#����.4`�Tb�MM��Lk����+6_�/`�/]4>���\���T�Z弜�|!�F���~S�5�S��^O�p4�C}������K^Jn��/bś����� lMl$���A�Å��ʻK��x�`�I�c�%\�.��2��Lv���>�D�A]z�B9!�UE�v�*����i�y)jL<0A�~|ZW}��s�>d5C�DC]�=-���m��o�1lu
%�w �����k���22oEud��C�T{�
ɖ��L�4
���#�'���@ϴ�-q�ci��Tux��|��U�ޮ���Q�R�l�{3�kE�7��  1�IQ��{?2ȭ(#f���B�"Q<t�`ނWSs�&�sJ9�G��۹�l�i��L�r���w����s�f��?� ��̉��X����/���V�,��GGOst�@�I���*v�M��q��rz�9��[�p4Ji�h��wK����"��jJ��!�wR�6G��L���l	'�nI@�1A�Uwu��Te�BB3�ec�{�����o�
�ΩQ���J���I�|Ę�L}~�v��_*�O�@���ޢT$�6��J���.���	��B�,8�|�M�"�(���E��փ�����d[��`��]�Kn��;]�����)=�m�9i�Єl�+iwSe��CұĹ�L}���m���M�q̬�Y���l�lS�������fM�Y�7)��+@vĴM@`�}� z����k(ϥ��x��3Qo��R����U������?ޜ���Zc�)���/��D��nZu1s/�o�!���C����7�2u6T�ҋ�b�����2��j�x��,�^��@#u�p������]��tR�G�8����'g�ʐj�S2A"����E�	�1s�����tss�?�i�ɍcuJ�m@�qf�Y�p�ߡ��rː}|~6M�FUC��b����D�Փ��k��+5�X�)�gd�A�O�q/�
rˠ��ae'��&2T��d��tdb�|/aw��{j�<F�@+��`mz�*˽j�����#�����5��lW�'��zodX�����L��"<���?=ed����ͷ?'| ?���B����b�¢s�7���Z�� L��H��ų��S��WrUy�1�a5�IY����`Z�����
�2Qi
4J(t��g�}�>H�"���;^�hvA��Ӿ`��V IP���5�*G�\��'�c�u�X2�^��Dj�������$��eL���E��dP�we�[�l�8����."l��&��z%�����k���h�^����Y�v������׋[�b��ڃ3~п�fV�[�=ܳ��zܶ��<x-��'j��2㴽�K��PkS>OR	4L<�,'�rzh70�Ex��%%U���!���Ҍ@� 1ߏ��>��z��W�C���~�Oа�!Db��~��SL9?�7<��wb�T��4�u�zo�V᝕�#�\�mr��@����['���f�cěU����U��	[�5��=�i9h?M|.�b�=1��'�9�(�p�˩�m����� �-ƅO'�=aH(�������ŴӬL\�PԽ����u0E6,��xu���0q��R3q������Q㡃��Q6�{nx�<R�"���	hmLk=P�����xO6� ��V�/��_�&������&���2�ߙȣ��;�BXO�~dGq�AK`*��t�6{n�!^�d�P�)u����SM��B����y�PC��lq@� �L��7�ʎ=�5 r�#�:�]��t���ߎ<�o�:�Top�x&�X�/��,�6�I������ ��%����eg��Q.�
�e��6�Zݬތ&MN^���S��ᓈ���]�䏰�Mb�W�3/P[/��9l��D���|h�:ϢEU�)E�+WE������{��Y��uQ�_���B]<c�1�ɮ��)���/J�↍'�/���b �`�Z��-#q��N�d2c���%f�W, ��ԧ$WHU��llݬ��Uqx�@c6�� �� �LR�?V����*w{��s��-��~~���6�������⩆B?�lM��;qf���@q���ML�"�Q&"R�$2Q��"K�x�~�k4k�(�#+Z�N;Q��V�d��.�LEn�aw��T�:��['2~L8l6�O�pn�i����
_��]�7��RC�`[?���uI �];/��G � 9U�͠s�۩A@ơEK1:�8-��������R,Z3��C�̥yY�);Ak��V�*��;C��K��(���f��#o/v�N�x���+�F�x��[_c{�3[Ui��s�$�y�l�$}�+���.;8��6b�&��@^y�AV��S�$����!~a� �&�����Q�?oz��V��'�V��d@�Yg���v�A�Si9�	D1ϻ�
&ﳷ�	d]�2�� �Z7JV�4�����wֲ��j�%a��2#�B��Z�%�t��c�]qa�eE�S{�ȉ[�CA�~��s�1f��hm L>�P1�A�i���(��[Ư� ��ȳ^K�ֈM�	�<l&�����"���akӨN�(�Έ��P�K��F���8$��w;<sp�P��<Qюܤ�����h��$�,mw^3�&��	�ڭ���d��e9��23�[O�u���Ut1�>��N�N~���܇�y�P C��ޫ�,���H-0�~^0&��˓J}�oe�+��*��I)Y�{��:L��:�{O"�@��e~�L�i��A�Y\�n���p\��E�����_����j1U*vS����=ж��mR�؊���@���a�=&B?�x�Rug�vo*��MXl�M�#��I�aم��I�ο���������o��P���] 0��rj�H��xʡ=����
(�ϒ�ā�k"����Q����U�8	E�#Qe<���Gθ��������x���f+}�&�oX	�/��_�[7�	�x�oW�Q�~ ��W��E�> ��Ʌ����+��ۻt�j�w�K�Hu_ڽQgN�R/?)�c���,��uM�2�x?[����PMQOX���&2Ǭ��g�o�:388�>ř8�E�z�&ɟ�^O>V�#���B`���s�hu�T$����)��x-T]>�Xi�T;%�� ����-6�[��k���G�v}�5��rс�t'�Ԛ3��i�X�gk�e��+�VP#@�(ú�U��Y~j3�6�*�X,;�X�X��,֌�'�Á������=O�K��G�a:%|_R�,��d�T��񅦓������+{Z��1��;e4�s��q�W\����K����)�d,��[)�n~�2e#�qxP��+��>�'�ރ�MWr�V�ir��޶re���n�*"x7wCUs6����粅5��/�`��?s$��i�R��Pbі4����������>un�;�b_�2��SZ�3�_��&�ֶ?����:{��T�����U{E
��7��-���;�`�?_r�m��B�|b���ͣ��ɍ�u��FЄ�f��'}��e���E�p�æ�E<)��=�%�҉���Y�����X �S��8mo���=�ݐ:�}�WY�0�<���>�<nh�Ƹ�J�(,VH=4�S�
�6���|���o�d�����&����W�)�_�T��i�iI֍�r�����!���8F$Vm�N7�R�m�j��л��M�_����ݞ���}] t��E��I~jGj��(v$�1'���y&I�b�B�ld���CB�H'X������a�ԛ&SW�����C���ū	���v�y�ܭ�D��)$�~�@ڛZ7�>ԛ	3���2���
uy�!~N�#;]�(J�Ƽ���L$26�es,���@��d��� zԂ&��鵐;���ϛ�\���7B�7���1*��j��S�v	�?A@�4���v�Q�����o�1�Vw��1���.�v2�q�+�iG�}�G���f${X*ڤ���Ck(������ž<a�MA߯��א(S9
T02F�׍�2��SƱ����j���=:u���q7��)����O�Ŋ�:��ڴP�Nszg�@f��i�(�dԆ��ػP����`-�u^#�g����������v�f�H<K�o��lf!����9 -yE��F�dV����k-�O�A�d��V�h�C�R�e�7"I��"e�~+�!#ύ0����h��+h�3�ת<b������?P�`�&�S֮/PT~OG=�Z��L٧<E�R����ϴ�T��_�:�0�X����E2�Z��e��}��	'U���|�� ��!�?�C�r����0��L/ ���+�D�Tm�<Xhc��zm�EYm+6�QI��~	�#��u�*�	��� �|(U�O��W�u�^K�������������\Bf7��\R�T�- �'����UG�Q�(ժr�wK��5��:ӫ��$YOE�������Ҷ��&c���#�Y,�Lѫ��^����B�k����a���wʟ� "�J������}D�\�Ϳ� ��.+�7+�]��0Y��#���R�p���}�1���#������/SQ"n�*R��stJ�:R��A�:D�H	��Mwa���m��S��BJ��s�wq���DF#���sj�i��N��4�$e�u����U��Az%� ��5�|8�asK ���k��VJ����շ�u�~?6u�2�.zŗ̓���n6��^���T�=�d�VÒ+:��<�QF����1���5�0b_etU��ݑ�{�\��ֱ]4����E��xExۆW <��ހW�E�I]�2f�:5��&xdQϷ�71�תe�G���#��GVD؃?@qM~��(8ީ�ڟ��h�����^�L�wz���S���6.���C��G;x�{�.#���[�+��/5�E��ܔ,E���9�~9+ҕ���P�[�C�ZR�#���.�A�;7uJs�@������Μ�P�Y�aFO���wP��i'��D��퉕�6a��8q1��4V ���������ae�(�%3��u7$��@�����P������ҭ�V�����V��f^sE�ezDZ�Y���x�M��'vo�؆E��{��<j�
���p�|'����y�h�!�O$�(u�<c2)�S�����^s�{�MWGƂ�e='�Vm�0i�{�_F�垶0p ��<K.=��:߽ļP9���U���dh)[�B�`.� ��xq��V����5_�շ�H3�iP�S)���Sk���h�����=8c#p�,c�~*Q|��)wV[�H���C��C�ͧK=D�U�}�iX<0�$�gK1�I]Y�J<�87�k/��^훳(��a���]�0�~���B��Wf��9�E=�@o����U|�Ct��Z�'u&"�u���dT�	���dR�A�՚�Ż���@����'�~81�h�S5���>���-�ҭq�I��vR�R���ط?c'��(ݭ������c��Nz
%����D������JhF�I�ƶ	�kC�"H��9o2��%x\�����*Y6�(��\�jAig}"*���O�x�ySD�p�an��ڦ���p'�.(��� �(�����'~��eP��U���M��69�[{X�긳�����U�=����a5p9*U0��e����`��G����d�'>C��f ��'�r�e�a�5@�i۵�sma>g�6-�>�S��R���z�]?b�Ta�v� �g�/��PZN�+(�m%�g@�_A׫�|�yu hu�(��Q�,.�z/�&F��*_k��o�r�����4�y ?��g��J}R�2��Q�$F&�	_u�m��-�)W�	�؊!���~�Ɏ����_^F�jFa��VD��ɀ�1��G��\՞�L��C��e��ߔZ����k�v8�4�Y'�DP�ARGQf���}e��zH���K���2�{��˂�x���?0{��囒F����[R�<�ك�_��z�IL6r]?�ذ�~��g�j���eY�rF�_-휨,��vArg
Y�%�
5�ؚ�t�y���*�Ȃ���<!��MT��%-_x�<,/̮�t@S��R�e�1U�h�^�=�"}�@�j� ��=��N�e�h�Iҗ囑�ݚ�˾��r�Vۡ��'6~�t��ja��D3����:<r�js��X^�Oz�o��<ٙ�)�A`5u��Q\&*��&�T@�2���׺ȡ0�9cr���!)�(&l��u���0c��"�=q3�$+���_��h
���8�yD��/k�l~;wXӺ4�a�Q��Q-k������'X�J���-=��� щW���	car��l�KؼS|�d���Q.����6@J^-���y$�~�� (<��3h�Y�d��2+&�xi:��k����f5�]|8D}m�긵�
Eq:�q�|/-Sxu�f~�P�(�f�]��Z5+�0�PY�*��0X�O���ˎ�-�~�����]�z�`����bT.�.8��Y��I������N���>s����V�E(��ږ��Eo����@"��g��ܲ�_�\o��(�2�ӻ4�Jq (�`-��3���N��&Q�8�N*A������0��t��'�{b���7�c��ć�T��v|�3��hйja���=[V����wL�C�s�@�~3c���1{�+�#�Q�U�I�-�Jj��,7��oq��q��H�o<a�><���s��[�82-6�0�/�JaL�o>JR�ua;K����S������f* p͸�]Xm|�'ZM��@���;�0/�l#�y��%YbeOO<l2��ލ���8�O��$^%F8��8�߼�U*O�8�d
5���=5ҍ8�󖤯���՘��R��\"�9�|Eϰ��d�>�J����K|`˫pTc���'<��	��!(����O**��#�ש�uP�*��Fj\o"�.2���s~g���Qs\���X�L��6E�V_�gL��x�~]|�V�v��*^y[�+^��9C�+�r/�T�){ME�BG!�$��r�,!cXh��6�dn f�T%��.Q*R����v͑Ё��tk�e�Z���Gr2�W�ː�E��|s(9�� ��R�d#��&6N�
� �G�l3�/1QUl��N�y� ��BŖ��P�5x[+O��'T>����#:#���㲅.,��+Q�"^g������z�M�����h����h*��27D �Ȍ�rr�j�L��:m�0Ŭ�|<�a�+����Z_d��v*��q§fKT0�6�U9QWж%���~@��Q��饸u> 6|�A|�`�1D+<�<�8ޟ�Q��L������}Z�̬��������R]u�`�ML�X��0O)��h_�c�VR꭫hʳX��&��r�ǥ
mI8&u�������"d$6k��oG���Z@�@%m3%O���ל�sL�@���)T�ΜHaĺ췺kB��xC�o�!�	y���2j�F��[��af*���5~�[�b��x�-U�r�#�t1|�D�hA���/��(6>~,~����b�,�Q`������B#��5�g�Xm�g��΀	��`�Qϐ
�R�s�޴(f��Ƅ9]%���EH���E6s?D,�6� �"%�H���daN�+�Q�)�=�:�"aa���}}c!�v.R���i�	�ڐ&�
����7�M�4V�JN\���$��ٌ�1!�rf�*_���gw��*�	���8Ru@j~sr�;I�Q$H�.��8����Ġ�N��V�~��H+i��`|�,��x�}T2
�,���:BT,[?4Rso��P>�d���'|�����Cl�����>S~-��Ip	��B]�/����W��9��v�%���ʜ��e�c>��,s<��UK��V8�T�vW�EE����ּ����:7�	��q�����~���c���}�Y�n+ϰ[ډ�P����We>әl`�Z�뙴p�o)��⪂�쀟�<�R�l�~�lED�}�	޹M-6r���+�����_�Q�NN����C �6IN�3�b�.`�#^���<���k��-�x@	TC��k'����A���^\����o��� �I��W.�y�`�����Im/N�.�Av�*`��:��e�_q�q�P����ҟmS�=(�mb��DǃWc��@��Y͉��]�ν0KY� ���D�'>tv7!��9�s�~�#�D��H����ى��~��ةs�� ��	4�Q푶z�]yP�"�.$6���� |�iPՏI�O`�*=�~y��q.v�뜚O&�\��SM�`I��o�)e�oj�:
��R����p3F��sƑ4/���y�w��X�|�~��ກ��,")]Z.|�YH�ۡ�Hd�($]q�j3�?��
k��I��0��'���$����L~b"��y��.O;�.դ]����NǬ�������E����,���!4�va��2��O��/��C��:܁VB�h?�ha+���YHv���U��il�C�n�	��R��ͷ���2KW{ȭ4!z/}��EF�a�@)	�<�.:��?�Q��hh1N��4ɏX!-�K�n�ߔ��8���Q���l]�e6'�'���ߐ��?΢L��̤���1R������c�d��P�9}oK��ǫ�o��a�U�߶�&��Fw�ȹ[�{�a�i׼�3��Q��mGh�}2�W8օ1rN�ܹWvľ��y�+��h�𘢆ܘ|��S(<>��*R� ��2���T����OKK�Ϻa�^�5���{Ѐ���^@�o{�j�,+���jil����8^���.{1?�e�9�Z�r����U������ť�z��|pL,Y9����x{#F+��9��D?L�.&�%�bd�2'�}��:��wl�8����H6����e3�8��j�,=/� �	�q�E�25�n�T�_!H�0  (��ޛ���p��G�l����z� ��x؋��$����z���K��a��z�2���턤���'�x$��c
�g۔���$Z���׊�e�vN�f��Y���@�L�\r�n7 ����7~���Um�]=v�f����MιmXcu�O�댔r�Y_�4G<��h�L86�P��gS��f9�^���O�t�1+��{ƲMa�;:���\ڜ�'[�$axMv  �E(M�Zթ'��h���E��6�X��~ݬ�p�0+L̓{�w'�j��������ѕ2��B5��ǝf٦o�V��+�⹅Lǽ
�FGo#�\��Or���iמ3����4�3�	�|��I	�M�@I��U!�a))�ϲ
e[IEM؏fD�g� ��iV�B�T�� �y�9�x}�� v`�Ym�p쭉x�f��LIp�	�]��,C��%�~=���*�Ϛ�˖����6[~�!R��u��I���R6�L9�:��. ��-�d���h�?6\K݊�L�5`��3�;��=� �e�1��D6ѲWB�/E	'x-O��1��L��6d����7��P]XC{���%�������A�d(Q"��D��fs�f\�X�S���:�.�׸J�U���0_�q�ʀG0w���9zh���l�X�7��}��0rpY.ռ��NHƃJI�B];�	�~�N�i���L����
3�����*�\��>#��_����ꆲ�讝�vӺ��lt����/1���+ȻM��dT�n,��u���ڡ�+#���E�|`�7��@���N?���h\c����&���j�w��Exڄn�g~S��>?�V�~�����r�)�?�����B=�/I��Ri ��h~�jee�fK��#��nw7�W��ώ��h�S1��R}+J͌���H%�l�]'�q�dͫ���]�!<�t�$6v�m�R��D�"��[0���[H�Hӥf#���.�&���ph@����$����T��6&&��SDc���h��-����ݢ�� L�KY���b7Iǵ�=Q��d6�W�.*B0��_B5xM���S�+-�a�Q�hI�a�?%�2�R�<�2�i;���p;8��FΣQ���m��E�_'/���xZw��O��L:@'��?M���9�<��#�;;���Z^Mf���-��V�Mk����J-Ȯ�T��~�KDf>�����(��Ũ��:?���Y�@�鑌�@��e��;��+_2R����i��Hb���ܖ�K����P�n^���[
�'�ɣ��pJ��ČCpv��ʚ�m^�N����)L?�ǳ�a��M�*���exk�{oV����sۄ��7�	�e'ɇj�ƞ��/���-y�=9f�s�`��IW��?�>�`*��U����~;�������F����΍��0j���3/��PI]�:���q��#PK��Yu�hkO ��.�-��0ti��E-��g���>��v'���dN��&�a߲M<�H��_�j�H��n����)`��9-�c��
C�1�w_�'>v$�i�gR���ɵd��p'*X��ϯKq�9���	j�d��]�����o�M��SY#@t��w�yUb�X��ay|uYP��o+�]���v3C��xH�bH&.�"�JZ��bQnAHt��`c٣Y�D���)f[D���G��b������a��qn||GV>�+o�N��j������0�ʼ�ѭ���z�4q���GM�t\���\�Ed�%�T/
\�W�/�1�h�Pz6�U��dX%K�.rvah�(�fΪ�/���)���| ��q��1C�Dȯ�r(&��@qXJ��T��@�j��>D����*�����-^����^X<�d�0���`���h|aI�8��/$����Ȳ�D��6*�u*wC�����Ɖ�pV��G���]�Y5�'��'���ߺ�	0��;I l����|�.v�#��3`�����f�R�P�2�����(�O���k�7�phMXp�/p�����r�ZHº��Ոx�T:�xj���v��#�0�c{i#� ?+��yؒ4�f��*�X_y�B�4�+q�P;�=ar��l�d�xv���UI]nfoz�MU���>�#s�t��@�i-�+�U�
Kp.d.O��t/{؇�nN�:�8�h���$�V)ld���{g]�F��|�+��\�zP�)<�GL�����"����s�=��?��F�8A��U7���=Y�K���=F%���9���
��\WrZnS��F�#C�7Qk&qWhX5�e$y�_�����Φ�a9Խ���)�BI����E�L���%���z��� ����ࣃ
@=�i���N�7�v6 t�y��Xw�MNu9<d�+{��2��s���|Chw 1r͟ܝ\�����n�/Mb>
`�H��T���j�2PI�zf�M�����;�S&eU��ߋlj�3bgi`�#�ic(M41�������(Ue���0�|[a�T�5MN�+�B��֠̍ǂ�o���Z�t6��F/=諵�����]]8����� ���10:�p��g�=m�� !��F� $��	������
?I�h�I����Z��*$b<y4�cA�H�6�~\�~�v9�>�����Qo�Y�_7�)��d���/�{�1`�Ѯ��\�a�%�M�xl���?��Ȁ~�%!<��^�T�>�٪{�WX��!��#W)�ZCY�k�V+	���A�bVE����j������Ka�lUXƂ��wB�#f���^7�A&eH����}W�)yJ�,�۸���z��G��Z׶%j����S(��,���HS�1*�t͌��Z����T�?�wJ�`[���{HgF��/*�i0�q���=�������Q	���CE���B�d�u� ,:�[�~� v
'�����JO�JDY�CĈ]d�F6K��#��iK���h�ۄvGi�Q�@F�o5=�|0�t �w�U[6�u�����}�y�x�)7_�F�)��8��W&D�R��G *G%V�M�YA��������_d~ ��A`��&�.���(��2$�?�m�E��=��]���=�'�F��Ў^��%�����Q� ,K���=v^(�oA^��k�ڇ�y*�	Y�v4�6��|T�TASó�]��'�Q!��U��������^x�vw*S���P,��Uc`F��8�ƪ��/��d��������a�f�v��w���?�$ M6 �aķff��z�B:8�_s�n'��D$�u;�f��c�#C���g!E��
��)�0��
��x�X����.��O�a#%��?F�m�Jb�(BK�J���ȇL��FFry�k!���
��iU�)���@���oj��L��>��-ȓ�٧o$d���`e4���V�x~V\ A6��l�$�0�p8p�!��ç|}�l�A+-$Ɂ>��c�|Ũ9�V.3ui}��|�!�egl�\�FY�1�WZ��5�}��
�F��G�ք�@�5bI��_/�zu�΋���4:8e+27 4Y����#=�L��g���� ���}����*GO��@�/��ҿ�Y����%Ҧ3��R;N씛��f�֪7ۅ��n��m�� U `X�'�h|���@)�
�f��/
r�;P��X;c}�Gr%�rY����)��*s2^�dS�C4�J3�n��"=Ѷ���[��w0q�kg9���Ɲ�!��%K�H��T"&%P^g%60�ō�J�W�X�cZ�o$��S�s�5���M(\�
�_+�%�*N�ȟ���0!]8Ȟ�J$��G��?t=�~Xo�z�aAr���� ��G�Zb�=hw��^x����Y���2�z��?S�И�D�[�H�uRC��x� y5J�* ���j�u����G�r2�NM�>A�l�Ȇ�5<��'���ߝ��ލ��g]�Ј����mz%Y��5�g�BK�[��i�E۩nΏh��I|N^�S�.~w#Ӷ���κ"���E�����r��Ϧ�T�Kt��s%?;��k�V��Iۏz�>g��PYB:p�[ȅ\먋1�V�u�l0A�u�t�g������n?�Ƌ��6�a�����������
������ŦE�7L�N'�	��ǹ�zr�<�g���Ac�ь	�|�g��J��l�%��`0��C¤dW͂�Y�+���ߤ�����#��Hn^�AwT%l�X�ԁ���-����ϻ�ŗ�Ij��a���>a���5u���N���ƁÜb��"ĆB�}3:���j�?��}HkYP���}�邺~���lY��$k:�I����b�:"2��DM�X�e�N"=�K�@lB݅��#̭ؔ��P�V��T��!����e�:HĿ;N���x��c�:�8�}���+s&bOǗ���I���	.q�tw'k�2����_j+sBC$��˲��3ۚݽڅ��HU�o��7T���S ��͇�U����긔���3���ZF8�^߄���q�0�/������bl�lRt��L�dnr�Z��¿�X�AW�yyh����~��
n�r��ڐ��]��f�.w�=�ۅ�-�)�!r�����s	aQڕ�mO����>��CCݚ �%�Cs�\��T@��e�T:Й��7�ؤ��͟A�q�\-C�C� r���#��<O��h�6|F�>2�P�������W���j��>'7�����5�f҅4*EWJ§Z<\�����ð1�f�������r����A�*�2�pQ֥Y:�;[խ~���!0U�JK��jg��{��@�Т���p�J�U&���sTU�����©j��{L.��]6�G;���>א� >�`�B��L��Fdq�6z�@�}��3�����mL�K�k���5˓��Z=J�k}�*���o�������$�x+\�>�Q��S>�9d�b�1�9��2%]��|����'0�	�3���wg��n��b�w�ɑ��4J�� ���O#�i��\�#+�T%'���'���4|���P��-SN��<����[GJ���ǂ�eG5#�?���fwʤ�Q��.e�2�&S�|�������0ճȞ(��.I�*7�C9x�>9D��C�k���K 9oV(p�vS��Y�c��2<a?/��^/#7}Bg�'�%k�r���&�d� @�,�8�r7�j bO�~��g/J=l��u'r�%Ԃs��HN6&)溊f�%��J�Wd�|��� �]�y,X�!��,��d���G�t!S�8w�t,;έG5�@
��&̈́n��D�f�w񹃅ɻ��d��q>fI�F���v����y��\g�Z+��3	�Qm��	�E~9�^(d�P
|��*�	�R���R�yY��3���G�R�� D�uQ�vH�o@��_*ӏ	-�m��t��`���Z��"�WUX�.ݘ8G��_]8�B,|�X���ū7L�o~���nw�8�1I�z��6���Ǔ�	O�.߇��q���N�y��?������ⴭP�+*�9���Ɩ��a)�u��yć���u��VV��`�>g���[ز&�;�6�i�)S	�A�Ԑ.��uW:H��O���4`�Q���h
��UUMf̥J2�d��d���P�۰�}��B�K�%= ����\�gǓ�.��ө�����G��ҶWt��������D�D,��ʪ�ʰ��46�U-b��Uґ]�4���_x�H��]�#���'�ϯr���:��փZ#{�[�Myh ���ѨE-3�1ղ ��~����]'��o,�S?N�2�Ϸ+Ӣ�����#+��)Q�h"�K�k�Z��i�3�5;O�A�ȧ��<��I�[I�X����ay<�V\Qu8�^����/��C2��^��\
Iu��"o7=��Y1 ���vԿQ ��9���^L}#E�ԅ�1�P���J#C�䄜����ﯗj���"�=��t��]��TW�!V�ԋ�V0K���R�p �ơ����B��a.�_ !���Yk��H�X̝�n���ꗇ�U�.�U�9���0��@��B�~�c�9!qr���9^�Z>��^sk��}�54Xj��U] ����:H$�
_��"+�ɦ��qE�r��c��O�H)bU^l���$g�;��o�b=0Z�#���PG�"��H2�q	�P:��o�R����x=bޕ�B�T���H�}CU����x3$XH�㧘S�v�����y|z���=�~�d��
A�`ؗ���� ֧=�}p��]��>��Ʉ����ٹ���#M�����N{�c��/ʹr~���Nf;�\�5����#��G�3dV�g����s<PMV�P��On6%�3.-�AP�/�pj/�\Tf$��Hu{f���d�xꁰJŰHQ=�X�-(m����)�yN��0�g�$�8�44�J�ʷK�M�*��B"���0),��9����$�-��1?��ԇ��3�̯�β����G���t�����͙W��.}�[߭�9�2��t,4{��$��W�������N	��X��O/|8m���a�k�!s��:�ID䩈L0}�/ ��E��y6�磦�r��U�h1�2�W#��3P�h͕���_)밶b��z/�*d���R��Z7�'@ۋ]Ӏ`=PeAv�}]�U�}!/H��I#�Ęx�$���R�9)���d~�3c�����Ɏ�W���f��Y�#����˄��1��M���9����%�M'�Z!z�A�u>����PH�X�# �>�Zk��,�d�"�~�"+<q�h�Ǡvھ�q�$���缴��p��|�4��i�![,fr5ɉ�S#-��Ә���i#a{R��v	�kq~Z]��q�:�y��-ݨciЪ��DF��yÕ�۫�J5���F/�^��h]�-��U���#�6xo|�=��EI�7�=,�T�T�umc�7�&��u�M�[��z ���מ�k����YSz�;�q[�_��6i� {�:���,O,�{|9*�y7H,f�_*�-���d�M�]���[]rY�tN�^�*���9�I�j0H��\BZ�e� nm}9Rx2c�����R�o%r^#	I�@u�ق��F�vL�.\�؞�w��y�<�+Di:�~=d���۪��OǗA���x�
��VPU�>�%# o�w�*�k��/&Ϛ��Uq�-7���6s-��<l?氨T"������E��$�s��E,��a����*)pf�z?վ�Wn|9��"Nᖄ�@#}=a��iDU52܄��Y��|��n��?��f'0��g��n���6����o�6�%�e�AA�O�T!E��X�k �` ��������w6$z ^�.0@~�X����<�Ih�M&��]�z^��,x\�M"�>Q�*P�_[�=��8�����W�����d�s�"@\}b* �p��;�r��HH���r�)��_WK&M�Ⱦ�{mصl1���4x�I�J�ok�tp�O=�Ѩ�za��"�L�7
T�Q�����n9c�+����QD�[,� �,'A:0��du�W[�*	�~(�׬�p�U�b1V�Ȝ��bT^>^Eϗ?1�K���Q9�!�31���K�ʟ��Ћ�Kg�� �5�����5�jGC��M!��Ã��V >J�W̩��8�4VXm��z�
~!#�]�C��G.U������	��9�j#EUr��Cl�^3���V&�-_�<��p/�{���7��7��5a�+ȅw��Fzy�A^D���o�u�$����d�k:Pd"��xk*#��4Z��S0�*�Ƿ��_y��Yq��}�^ն��iѢzM���*��?�{��)�yW�"��Bw�"s7ņ��S[u�Y`�,���*km��1%�oo3%���"��޺9f&�/�l7VbWVn������{�Z��[�v�z�h�)R
h���2"�}����*�O�M��t��k�y�g��YF��]`�����(��j��"q�D*sd{r��N��-��!ӥ�Vm��m�P��ױ������%�;�XjaB��[�ycڝK�`�@ �'hbG٭J4���]O����0��6 ��\�ve~��y#�������3��Yl��Ozٽ##��׏���C�Yj��������ͭD��|	�­T�G���TڪmGǖa���2;���i���M>�'�>p�[�$��h0I�Ɠ�g����Xt���UE3�h&�f�?��O�\KB�qS� �7��h0o좌+��֔8�#wT����ô����_�6��̓P �ڿ<�=җ���tN�2.l�^��L<iĔa皙�0!:ۑ]cz��:u�rܻ_�W\3wW9!���4���2;<��D�_Y��y����Q�1_�B�֖'����Ct���/�*R����QY�?�ٶ({�P�p���ot0�0��J�mm�J#V)��ծ����5��4q��7r�Q_aسΠ9��8�D/+� �#FȃO������P"FC�a�JU�iU�N��<|�4?����k�@�&��1s�I�ɦVNT
�s4�^T�H��J��1Yb��sn��"4?d.�ٖԴaTQ���9�F���})F�8�9���2��9g--}��Aͽ6M�[���D t4�i��rX�c�c��r����7ୄ��]�}%������W$ڹzԾS�|��E'��FE��9B}��䥮����i�b�r���c��˦(��xyh�!=�������*��4A���' �e��4�.H��X6��&�/[�g�".�-�m��U1��!��?��cҠ��?�l�� �����ZL��Ė;f�_�W*��V�b��`�r�{8.y>ݵi����^k�4��E3�|%�,��ҨY�(~����������yw�t�ţLzF�E�>z�7z�3q� I>�?��5�!�Ě������J��3�su�s|�!�����Y��w�7�I#�PT6���If!691�wz�&�nm1�ʁ���
n��ZL�<2��cߴ��F��2MX�
��Ƒ��T�}�y�/2��,�b������f�av��Tx,�˻a�PW���w��ïڙF�\�0�
�rrV�
��h�(7�f��^�u� ��[�.QX�:2����*�tU�ZR��Y��T�9�8KOW�;Qޜ�<p�T���X��D�e�X4�z��`��I� YM4�E��C_"6`'�CV�D��it�[/'T�9)�z����
�sn�g�ŋf�����N��(��}�n+�Et��=�DF�����o�AR���/Cٚ:?��ɶ�@��Huj����$�_^�r@�1pZ��bk:��ɭ�ط��E���{� &�] iF�2;��Ū�D�>�-V�%�v�|2��A3Y=&l�ꔀ0�&p19$C�	��c��R{�p�
����P:䊭�m��,,ms��>BZ B�C?�7h�-�p:=H8v��;?�)�͝�9�c`����!B
�x�d�`����gE�`D5^-���>l���g*����6��B����<G�ML�wh�5.I�����	
�����f,�F$��QL})�9m��_����z����j:C�?Wo>\�*˕�z�����p�܇�V��op7 Z���AL��w�~��9pNI�,�Y�X����,+ 	����o���D����0�R�":$5&�ۂ����6@�h����{y���R��?
*i[%_���+ZP+�õ��%�Q��$+���c.^��fj�]#c���:�4 �,�=(Rh�4�(�	��2��R��[��v/��k��dJp�.=9��E����135�x��v�0Ƨ[��B�Ƨ��5�Y�{����#*}�"^uՆ^��D("�ն/d[()��K�j`����o�`�S<I�Y�w�֖_/�0�-�̅�E;ͬ�Ҏ볫s�qO�v�)�̥ngn���t'{���tr:`���s�{�Ǫ��4w~������ -L`���v��(�5�`r�X����@�O*f������#,x�}��܎����q�lw�H�HX|ɣ��'��蕰Do�i�C��J
pT�CA@�����ܢ봘P�#��]@_�mqh��8�)�h^�V��w��P�g "��f�z�*��̮��s��Qh���6�T��ʐt�;n�hרN%r���p�'+�怂��v���p,��4b�%�K𹅒�0��;.�}�}>��V1��_�~��ӎ3���O޷_"w��S�YٲcfWQx�|�u�O�v�mQ�h#^�NS��9�b�m���:��5����{�:�F��?;E{'�^�r�V�ī��I/嶱�'�o��0�]���EEgo�2��ځ���PݪA�3�qݤ����!:��t���4h�w��!�oG����q�Q�1��y"�$�/�u~��N1���)H�r��H�]�u����`�q���Aچ4|��F�"<�O��
V��3�ڹa��Ь"^�/��&k�pk!iK�8��H�%�P�����OI�uW~\ON+*��Tl����zɨ!!ck�$nӖ�x��%��x~��g�-�\U�{�t���5�6�cy'pR�&��Ge_���|ۯ�2�c��_�����D-��Z��Gܚ�6�Ҽx�Xꪜ�|�+�qVC����Μb�9���!G�p���V�����/F�t��LBy8e��B,��D���&ߟij������Ţ��{C�\N`��IX 1�]6�r�#�%'P�U\�"J4{��	>�K��N��ݚ������~D���:y��	���Qs]}�0��! ��j�����F�M���2�n��.�5(DO����N��H��;�Az�/��y<;�c%���
)H�D�v"/��^���<����1F�~���7߈/�L #�_��̦!�Ϻ��T����U�ֶ=�@z�sCoܩ`_$8�N���_Ϋb���Hg�p���CMI����Xoq��kj1����Z4 �$`}R/��Ns	�"���M��l����`���2�S�=~�v�-����9��!����3H��4��U�� ���X2���(�"�Q��b@\hf�O��/�N�x�>��D#�!k���,�>@Ɯ�/�χT(aW@�� /ȅ�j�x.�,5�:���w���u�¯�U�^��ĔA�^^��a:(�4.���7�O���+-7��V�ĮP�k%�]Q?����Oe�^���F���9L�[sC@��l�l��HNb�Xʟ�����	�sw71�F@뼦S#�v�\�W;�#0�pfH�d��r�p�S �J�e���^�C��N�s�����G�1\j]����-���
��B�[d��
0P<���@�h!�B�Y��z�G�LE��[s0�jO��̶�]�h;[y��R���U�į_;�1$b��j�_�{J�|���00�_,�R@
��zБ��w�-�4o:�]U�矁��y[� DN��H�'k�;�3�8�C��r�*n��������)H��}�ӕh�d���50�����4�O3)	�_��T��x�6^�.����X�����lF+/x����@�5����/H�DZ�`/Mdjx��wBJ��a!��:ˬ	�d�	�
;��M�|a�-���^M�ٞKc~h��5���S��\p^nL��#���W�^X$��'A{�5�6�++�8�+0�,�M���V� �����G�ȘɱΨ�%9s��A����T��*�[c0G��|�3���$x�ц�7�lM̭;c��X���2�)&�4������RClB./��i��@�6�pZ��k�w�|+-��I��j;m����/�obc���h��n��<~��b)�4��Xgd�+��������%l9�Kj��	���oP�P��]����������Aދ�VΛ4��E�?��N�&|�U��|p/%���Y�$2N�^�z�,���F�E�=3j�L�z�z�s�_O�ODjV'g��Ė�	�n��	9�xG��Q�M���{�R�L`�-�n�V��b�56 �/�\ؽ3'ɱZ�5��Z� �6�ؒ6c�a�y�v�Xlg�MI�W8Y�� �{� v�~L��,����wLH�㬏 �KVq��3��Lx�1a�Q}��X4c�=>Fui;,1I�?�#ޅ��ܧ��E��C��uEeC3���n|ۦ����S���ԱkΥ�p�[^�ymo ���5;zi燩�{�_/��5|�p������d� .E����c�kdY@��t�'�3���u��A!��\E��^n����mpiY���q�'�J=��!�l�t�|d(E|G)S.2�ڔ���'D�/qfY#� ����+�7�RrL���]n<vn��i��+��2��9��3˽!˙�QpF����%Z3^5$��`�=(����y�"����ĳR]:�wD����!U����\̓�V��N�d�WN5H���Q0���#a�;�	�:,!{�.�T�P�+���.��Z�+�F����[C�Э*qO���L����	Ep� ���g%�J̘���'�{k���k_C�|d%��W?��6������@����owwn"�4��Vqل�g���6�V I!�M��Ct���/�!�Wv�j���=VCs[����M��؜�CS_���;���KBUD�pR���)��p1�Y���K)�I�zm粘�
��������C�q�<<	�'*v9j&
���,��$� O���������xBq��8|l͋=k\2d\@w�|h�Hmcƾ�qw?V��nZ'��"Y�iT3r�cÏ-���}�~���\q����:�ׇg����9RI��v�;�I������F1�Ůڪ�Խk���{{4����u��Zf���wf��.��`<�@%�!�i�]L��� �k
�Y��[}N�uY(غ�bu�b���>����8Y�^���'w�Qh�V _=����C-��:��T�Y�|����A>����+Jeמ=Y���g��4U�GY�C��m)O{LG���ޣ�=�j���Q�/�*�+�Z��,V���N�� kEnH�@�׻o]�`i��,��gn��H���r��	&po"�a��D�@���?B���
�yl[��S��?�����&d\k��O� �<�[�C_���c�]�f�U��7���X���ۊ��s.EӉ_E�Ƌ7�����u�w�ᦀ�*�&��V�����7��+�ӯJhW�j-q۫��f�|�
�p* �B�z"�Z�\1T���]��ֆ֬vHV���O�>)�*��m�u�$��l��u\�����xG�)K���QCl*xn��0�D����3�|�S�*G�FY�g���]ގ�^;؀k"�qň"
d���@`�Tm=��b�|�[��Ri�����DE���''@EpF�jempˉg~s4���d��+�]�s��_\�h/)�X'Rc}����������_�O��mZ�f���t���?C(?i��1���x]��jJ����<t�f3��/3EG�B�=���l@>�$	�:#��*�}t\遇�v�G
��V@z�$�� q��oÕK {�Ɓ*`��$�ɩ���N���}�fXx4�W&cz/G�=�D&�����%ڗ(MLTӜQ(�4�+���p$����\�V[�Q�AV��ip�5�|흫��*ȩ��u*��ȸ0ZL�����e�
f������h�-+�k@�u�8W7/����������>�6;����}�*m�<��Ż�V_|X��Y��
�p6,.ο-
�`N��͢йU.��U.5-+��N��2w�	N�"ӑh#n$D�˥5gAo��ׯh#�Us�iwS8$8S���ng`R7�Q�
ܻ��ȵB�X���u����8����'B�9t4���ġ��w\ΐ4�hqM$|Ert�>F+7���1`A��15�g�օ��d����5���%?Qʛ/��L譏$��紐MO]6kE��8XH{�BX�	�ȣCx�3�;�<\F�8�-'�ڵ�^�J>K����X<�5�� G��T��.J��Ԩ3L��S5���?n���8Q#�6���"��	�lY`p�љ�8딑��a���BP�آ-(-��oD��B^r��r�A�nЗ,�6e;��5��xE>��IZ^���/���y�j��R&a�Ur�U��p�n�������*�:��%�������P��&'�j�+�6�(�(�*�I���3W��������G 4�۳�\�U��}���>������!T(���^�xP:nb�CpL�S��.�C @��^��;��6b'C/�c��l�� .R�/��΁��B���"H��bwM�wF1��Z�t��jk\RWo[J�����	=��7��;���Xsc�0]qN�����Vv6Gaъdc#���+����W���;�\瑯���w��2Y�7�`��P�w�z�8��|��-ɑT�t�b8(u�q�����]U��I{�c?ʝՈr�qr%�a-7=�v/���~�+�p�e�E�w`��|�M�xߪ���[�p����7�E����Ę0Y���M�� _�ѱ5�+��	/���w��+U��H#���`S����JЧ,�����7/4�1p���{e�?����f'�	'3��[��:qEU1)[-�ϹNN�:\�6���ui�!a���@l%�����4<V�;�å��q���$(Ĉ7���@����d�g��G�%ɐ�F��w�k��"+��v�TՔ����Ś|m(���`dYSҎ�D��f�}�/�ʝ�1Rܨ��?ϳV� *A�jS:N۱iE��]�CXβ�Jb�S�yr���2\�2�T��dFTqם��	r���k$�J!�:����_C����>3"2����QwZ�o�����/�'�x^TCTe
k���{�:e�GOOiL�E�Jʿr�H>1�@덵{�,ec�n���J��P���bp&nZr�Ey��g;fIuml]����d����d��r��|jf{Q�!y�#`E'�\PB�bd:c����\�W�^S�T{t���YqҭX��$�_��>FR]�M���+��X�x�N��4�!�YKZ4�/�ћ�ˊ)�M�T��[�1wb��^�W!Ea~	��Cΐ�J�|oU8�.)��Y���#�4��:�]zV:��n�E�6���L�e�v[Brk��z��q��c,�ɏ:Z�`��S�}`��5���Q
�-�O�1�:�bq��u��U͙;�]�3VL|<�"O}�H �Pߛ���)Ӿ�rf����iU�����wv��c�r�_Y'@��C&>�k$Y_7�qsS�d6jb`��Ϳ�݁v�?M9��/1�CFQ=0�:&.n0�ý��oI"b��i@��a[��ʲ5�_����;E��BΡ��T��9�% ��淭]]�0\F"�bDH�����-va�lZy��-k(Q

�@aȈ��+��.kp[;��3���w�%'�ΝՉ@�c\-�Y D�k��-<H�u��l��N�� �5~̲HufE����
jmc�ZG�7��a=��p2���F��EHo�^-�v�ms�8۵�Y�I��Ĭ4�x�S�僣b7�x�V�)9�#1��ⱷ_�i�
�6�a~�A�QyNy�?��a?M�v����]P5�&�a�z|���^�8~q`o�T���c����Mk��$!���f��a�J���W�D���K1��m7�[�<���7�ɑ����n��*^>�ZX��^�&ʨ��9�Ѧ1��V����c��^;(c���v>1�vZ�[lc��R��-��6$:����$M���H�^c�������S	L4ey�k����$��9���<���=�W����l;��w��Xl������_a�G�a�nH����b=��>�6�ӂv{2��Q�ܖ��n��b�a&��-�n)�
q!$�e[� NBjvi�81_Ff^a���r�&��c�e/���h�n�:)�ʞ4Mҙ���
���t���^�z��.I��D��kwy���NQ��B�(h�(��Z�j���X̀:�s�yV
���㙕�V(,�A,�w~h>��-h���-�2�NR�������O��`x.���t��Κ�oi�,P�]�D2�:iq�R#jJu~y���k�<<2�l�a:j��p�bw�i醭ߤ��a��4E�	|LΩ�Ӳ�>;}lL,݁�����(�۹x8�a>�
��SARZ��a���aeu%�'?�O߻�s���u�=Z�!�W�֗�C�:�;�r=�_ZF_��\��_�y������j,X���ry�^�,��}��zӆa������!��7�Q�w�=,e29h�(�����D��}�62�����r.�Q,�2��p�a�-J��������Iz��6���'�D*�����ӿ��FΗ�"x�$��J<��Ti����e���֌ք�j�-��i�bk�A>� Qn��]߽xD��.��ŝ^"dI�M��mG
��mu���7�5��o�m⡳ գ~� �\�km�3�E��k�H�[�c����B(��i���v��ZT�=۟"U�"A�o�	҂n>H�
U�(��1�>����{��y�Ѡ \�<�����&aʂ�1��C�)�t|v+Y�s�alT�(�q8�Z7��Ji��q\�s�E!��=�G�� 	���uB�0�=�i�95j���;m��e�f���\!c�35a��S��!���VT��+�"��P�j��#_�U���_�|��\=�R�(5`N<M4���9���+t%T+7�%���Op};��m]���o��w'6�F�!�K۵�,�w���WP{|�"p����Ƽ���/�t��h�>o�ʣ
m�Pz�=8d7}3fu|�E/5I�{:���A�A��D8�c������qy�`��d!����t��+i��ܝ����m�z�*sl"����ޫ�(×�������+^[�\�4��@PY�'��d�p�"�����X���q�iҡ�/ӱ��$�zV�i�/���3	=����F	���9�/['"���GN�
���~�� s�F��0�\��,�	9J��/���vW�d��z�vaoA�@lH�k4�I/�s,��V�%�n��]���V\	 =\�ٝ�X6�zT�起�0+�V���h�U�uX�
��:�S�pN���;)�H$��=�h��n��沴�eF��$���2�)��n�X�&"9QC��v���X����8��c�E0�*v�zr�K��7y�j��=zx�L��]C��U�� t!�,�Fb��.� ����*�}�Y�0�H(w�J�b��7�H�8��M���*�k3F�1Sx�"��2����B��ۓ~�����ٝ#Ng�/�+�;��8�1�\tI:��آ�;��x��n�itʘ؍�ꫨ�]�����+Qv�i�od��rd��g��kϮ�ں5����ڇr���q�F�(�֒�\r-�,E5��ı��6���{Zzj��D�K��8ȗaf��)Gl_��v�����b��>#n�����wvPF��'�I.�����:��
krBg<+aB�ƪ/$R����׷J`���M�rq����~
��Q�8wk+�]�%W}��њJϿ�%<E��s��aK�j��'�0p�Gm�{h�֭#p��C.#e�~p����@dkYY݌C=���x8�j��}�4;9��Ū�ؠ@e-I]�X8��������V�6�xô�/�9�Hĺ=r6ݸ��TV��:��"���S��]2k���n����e(���%�c�/a��>����ԁv�e���r#���4gz:����zr�nF[rL�:q��P#F�����\6 �!S�u�g+	���p䆌c�\F^VM������@H
��<��vQ�h0Ѹ^ڡ���)�F{�BW:�rV���!��=BY�-F�p������i�%�z��~]]�Se$!v*7��x EۗD��޾�`�6�Y$*�;a$dMU
s�EA"��ɘ�7"si��U�2�7.̀��R�$KR���d��[묌��Mx���U� ��+0[^�+�:��h[�m���G���.X<}�L>��9�t����&/K��:�?%L�YE�0&�V�4E��AE����N��j�߈��/�軑:DO�1�q�\�ah/k3�[�:�ۨ�hL��#�ʴ��jy/�jr�IY���y.l�����ٺ-a!�w�,k:�:��A��1�����(��;-_��Bl}`P��?��p
0*ԙÏm&��!���[�a%�o�9�F�i0*�}u�1Y�$%��O���������'�h�������S�G�4��FD��n�g=���<�1��w@�����W�D�Jn�S���8���CE��a!	����\��Ao�������'��V�}r�S���լ�����'�i$U���!=4� (�E�~��#f�>2�1vM[� U}ٌ�鈎�i
~Q�x�BB~�G�BY);ߏ�	TW���{�5X�n�gM�2#	 �B�UZ;�dHf�;Z�Ҹ+Cm;� �o!'3G�,n��#�[����-�d��PX�q J�\����e+�ք��[�O�E�;J�wt�����gOPG��ӫ�k���V���.������sS�ha�:�zt8�@憽b�dx{5Щ?�����Vkʨ�S��	��a���P��Y�O�K�_�+CF��D�rf�sN����Zy����ATW?��H3��Ɂ�}?6��I��90�}�6�,���Ep��L�C͢�5i>q���b�����W�ɚT�ۋ(|r����.��p��� O��O��o2|̖�J��i6�w�!�!;0���ъ4 -no��s��M��;�mITD����b�q��{�Q5���`jJdlNj�w��SP�AZDԬǇ$�֫��j��왃�y�Pk�Y�Fli/�$���9C�r?-!K��i��Tj4o�62\��o��pQt�`���>}��ԍ���NGN��$!LT�מA���7H
	[�R�"?4Knz1N���l]Y��dd�P=?)��k#YR�ѴE?o��C6�+������{~�������c*4�G���T�ͽk�[J�J"�ڧ�g�Ouf���-a����hLKe�{~���K>�@oX��A�93����A���cc@G���$�q	�u3A�I:�s���H,�B��'���n|���'�U��ƒ�G�x�����<9�(��O�9y�s��Z�ȝ_8�v!��C�KU�3�S����"jbp�w���ju�\�*���X�_�Hh٪k�o�"���->��Eq�� �fl`w��ȭ�Wai��2�>)4���fKd~�5���r��<��u#]�(f�%G�c���p�jw5
"�;oW6#a��!�˗��*xE�@���{��J
8?����� �P*Ky�ۻb7����&�,@h"o�Hs.C�t�(�n�~?=P���,� �57(���:%�{A.�}��6%|sўOY��~x,��U�GͰ^h���&l�� ��oW����4.մ�#�Q@}���7"�����Lo��� �T�y� ;��k��:�u׍1�5b'W�:�\��'�F"����5�߃��a�Lz��,��|]�F�|3	k�� �g��Ӟ,��M��-�̂�q�s�Z-�,!�#��AE/!9/�_���P|��uT�1XZ*���)��B�7�����&�"_8�θ�����%+U�Aۺ��Q����f�Ot,A{�R1�Y�s��V8�����:�B����r�a�U�+f���Ɛ���%�A��;�\�W:�8%v�Nx�,I�sDtX�T�l����`)� f�Փy)#&���X�X��bg6�����2V�6�x��3��%���`��.CI�lw<p&A�ո�р���0���(�}�	�MGO8���
4��3Ş�5�]�f$H��->��r�T�@��dwN��P-�0Ư�u�%'�ô���^{��P�_��銒�z��9,�L�
ڏ�9fĉ�p�����.�(77�������O���X�������:2(�y����Y�s�[=,�tn�_g�\�TG�]�Ɛ�X��ȷ��%�	0.L!�9�K�s�����Ʈ��l@���do�*W	P�m�npO��]�=������9�/ǟ#�-mG�d�k���l�7ǲd�+��1�\�����o�~�M�P�]Ld��\���6G����H�ҒN"R��p�wqkfgˍ�p����[!D���<��߁�|B�X�Uq�g)�L���(�f�J GU��;�(t4�/т��R< �ջU��35���&�������Y@�|	d�Q�6��9�	�.$_�������/q�b�0�%�;�,�}O����tp�O�1<��$}��>HpB`���TM����h>��D ��V��#�s!��U�_\�^���|9���gd�8�� �3z����h}jk����9)[�.L��Y̸�d4���iKuX�2������~�l1�	���Fv����!�)u�g�N�W�+�G!Z����v�t�؄E��+�g~)��X��m�UY���@��R_�U��-{؜,\ �T}o�߃qˏ��ږ�PZq�Zn�:�j�18�|e?ZE��`�����1"�?ٴ�w���t8�E�3��@��w��O���{P�F��k�yȘ�1Bџ���Rl�`j��.���4�e�xA�K�O<��:��
O��ޚR��?_��X�Ev��<'ғ�OP{��)Ԋ@S�����6�2X�����H��9;bOR��Z-z��6��'��J��LJv�.��C��Į�K\C�3ɺqa+�/Q$���WѮ}{V�<���~�[���%��7Z���\"x�����pJ&�"����lVK�}{qrRv;��v���(�|�)QM=�j������;i��m�3���a�D8q�[V�<��Ƨ�Z-�������z2��v��LO�e�7����eZ�=`D�h��Y�SQ��Բ�Z��o%�ᑽB��9T�+ա�8��5��ԝha�d�7k����Ă:6ҡ��|�W�d{�j� �9|7B���-N�Ri�܄�x)K#�Q^O�8�S_�߹�v�ޟ�S"��ӂ��n5�t����+��|W�6p��¶i|�v}#�N�h}��&x1�7>�{=��Ǻ���	ŋ����%���IX'��I8����0ǯ��b�,����r}�A)��hҘ{o�gzyw��R8{#s���á��"'�C/��,�%�Ѓf�
��� �u�����ij���6�"}��~q�(�Z6׏{����@�d����v5��g+��(���A���Xa�mIBK�����A3�~��n�^��Oh�sH�W�]ϳ��{��:`:00���^
�4R��/kΤ�[�B�&�g5����	���&<6�4@��zo�~[��)�髇�ʎ8Qx%�ש�2,}�if�c�E}SP_y�n�ڃ%�=G�Ъ�ĕނ#�fL�9z@1JC�7�����EF߭��.�zmݬ������8��{
�-]�
6|��#�gf냷�Y��{rU�V�&�t֘����@%+�S�`xa�ƌ�������G�u�yzf��I��I��T$��S��Q$�A��͍��������9G�6���͒�v�4��v�\6�or�E*	�@�,c_NeW���#�,�b�bcg��Kv���ԯ���N+������Pu�)��.��ޣ��]LWc��,�7b	���DS�j'Da(���1��٬�������|�'�����U�D�QT�º��x=�<Du��Z�w�h1�J�F��NgR���	��j������7(lD���dW^&��>����I{�ni�����1�^D˫�uy[kg�a��K��nx/��b�G��~�c
[�q�t0�H��`�/���/ş��g�#Bt�����7QY`.�����L�;�]h�,̉�g:o]��	���T�ٞ?�����h��T@�+�;����g�`������]�/=ia�u	�!���������`�iC>��+N蘏��G+k1[��{�n�{�'�ݨ��ߴ�����MQ~Ivf�u���n태b���-;��,첑�~�X�#���̜�x%U�?@�&cGN.c�p����d��c�ϱ�	��D=������a��nՈ���]w���u�� ������i�(�K��8�Ǳ���$>u���)�w�����^	��;۞�@��Xl��YxQ�moYSx�Q�9X�z�ɍ�`�j�\Ri����5eKS���>��0l�w���W>ӕ���ؿMbӷ��txAb�>'r��G�1�goh
��,\�:���96�C
���PZ[�f?R6�wf���������+$M��P{%�+����e�Ί2xI�?�7�E �kRsZ(4)���<dڲ�!�����+�������T�ܿ�7�%ʉu73��^/��A�c�1��@|��_p�^�3��l�����E�C7O���|�9�_i�������i(�%pAgQʘl$6�G�;�f%���I��Y~���;5���z�I����c֗3�2������aF��� �(2]�m�Kz�[Ё<��u� �|��DP9��HJAʒ-�����9|��
��0�VL�����As���M *�䅙�ŅU�%Z������k� ������^����2��z��r!'X�cL&���{6�$�
�{��v>���U�<pO��,4�V�=��Gψa��Zy���ٳr��,���P�,LL���-i ��9k�-�t��>�	�;�=Q��^���И��,�g̲`�VG'oJ|¡�Թת*�����H�o���D	��;��(�LQ���5Ztt�Vi���f��A�%:�~��g�� �zV*�m?��߁^���b�-�jfQ���W�����E"�w�e��P�s�\;�Y�H����0����w�j���iμ�+E����Ge,�2Hi(��u\e������`����[���c���>�핱BF�>*�d��3I]�!(�X��ӃY<�r���;�'������7�o!_�wCއc &��K{�+Y��~p�Bx��{�Q��`�O)Q�N?ޓ�N�߭Y�eU��EX����7����������a&c�lz�U���t�"�Լ-x�_��pD�-?�A�A����)���5��<��)&�L�w��ʌ�	&�3e�Y��K�*Wv�v�7,����=߉L=��oe3;^��=K8����zC�YG(kc����JL��A�'M�!��Pֺ�45sh9Q�_>�J�7��Z� x���D.|5<@L�5��1�&9����;�NA>�	��&��[|��~�6'3/�M�p; �QO1x?*~�g�%��������x��*V{��#1���-3�e7G3UN�8��+���b�`_'��ԥl"�ђ�|�Cw��2I��c���P�yX^��<��<��Bj�������̵$a������KM��Z?�T�9�XRY	�ѯA�}y����c��(��pH��;ҹ���p�v�$���hp)�S���xuXKH�Mk�P�n��;e���q��
�W�rP�Q+�_qgKk�gL�h����ʢUوaA�!0�����ii"�4�8om��Q-��\Yt,�\()���fu��%�W�[���ė#jɱn��W`��J���>�`�=���f��:޶���z����C��V7�J�viTg#O�\��#:M��Wgdw�j,�s��!�n�Z�V9�U9Z��,�1�G�U�B�dG�3���9L.W��P� Va0q��H�����\R��!�+���9,����n�\��k\�7GK�@T�  ���6Lp�=�
�~��i�,NT��u��0V������/��?�U�1��hrT�"��$��w7B����<��0X� ?��n��ya��)&o�hc�/C}Wm����e�[l=:S;ǀW��k�u=1���qK��'�!9o�}�h����N�Ǽ��vu��'������̀i�(�71�dQ�UZ�X<�/�y���N��w�O-
�-/�퍲�\y6����i�μ�Z!�WOmd��8�ҍ�ul�+ݎ��ƒ�K�T��2)["˦�?>�;����XQ����G �hg�a�O	��-\@�*�x����t�,Bt]���!�U�V7F<��c`�K1
I������ȼ�(�����tF��#�mS^6��i@8<%�S�`5��mG�:��w���'��}o�҈ڷD]NzHC���LK�����
n=�(�b�82��.}�����,��T]�LD=0d9Ϯ�eʵ����yB;� Fٔ��n��E�
)l�	�y��=׽|0�c������ّj[�i��Gf@�qI@eT��gF��H��'���-�KV����Kr��gB�dU�e\0ET�bn��#T���54<��ZO/�w�����<B�r�qi�8�����M�+/�]fg?)����y����α��J0������ujp?�;t��S�X�2G��9-��z}ƤE���u�cK�x��6�foM�ny%C�W�̳6F���	�Øj8Q��u"KY��S��"b�/��?��0�A�s*�����,%T�HZ`����ו����و4�V���-]b&A9�k\�)�Gk�Y�JBE�p��^�-���^�.���������Ц�`Pe�q}M+Âf3�u1nk2�&+p�������h=�4cJM��芐C1�����l^�;��C����_��}Z�T�z����H&l�ן%�����v��gO|�h�]�ٓ+�|Y##x�D������5����*OZ���z����p�����2_�+gi�gH�Y����Zȅ�!)�`�jP�<�r@�]Z]F�ŷ�A��?ʛ_/�D��ᰩ���Obr�
Q��_J���"	(��!S��7����_��=N"o�w|���/%E��v�mҿȆ����6�����6�6vbK��