��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&Ű��=�b��vT6�4��L�b,	/,A��"⽰k��b�t�u�zU ���� /��QU�:�4l�Ӟ�l�) ��$�����6�Bͣ �%>����4�p�ayt�J��C�`MW�Wd��c���lҨ4�!X~��V`�]B��楂Y���H\(�2{�1A<n�9��g������(2|'�n��ݡ�r��l��e�O��9���S��nwA���@�*ں�Z�� jU��r~b7W��t]5��g����T�[�tdJy��Ğ�i�\�$wO nOp��C>DU�8S#~�
Xv݅��
�Q�`Q�dp�*A�X�P�zs����3�$W����n�dοUƺZkEϦ�dH�<���� ?F�S��|TT;z���H��q~�'��Lh��%Pa�m1]�2nW�H����	�E29<-���Y͗��>w�F_�:�W�u�����+t��^ �k���|��L��!Z��#N�h��E�v70eb_�b�8����<��xƽ���M8��Tbȣ�JQ�உ�r�2`}�{?=%
�#@4�|#�y�1��uz�&ZH�1��<�j&�X��-!)�,{J��I���L� ��Q�΍r-���jՠ10tSZ>��[%�{��4:�RΝdD�Q�Px{�E�Y)~z����Ywp-P��r�?� +&w6�Yh�g�^���
�F��mi��(�A�4�/%w�?a+����H��H#����8U��`]�^��Z�M~l�����ת����(����z݃ �O�D�%Db�Z��:�+}:�򰕿�mgL�D�̀u�`�[W%v��_Fs� ��Lz~��Z�.ܗ���
h����H�$N8�!(��ʼ���׿!  �I�����U�}p0E�ݡ��Щ�}�$�>Y��@�o��L����k���B�CQ�ߞv�@�%;1���P]|�	j=�.!*n�&��P�Y��Q�u"��Կ"��Ԇ����_�tܧ'DFն!���2�>��.["R��A*�!*.ȌKp{��c�rLiгG�<�� ��x�j��}�Z������^v_�Í��Cڷ������F+`o�+ohSh�n�����D�/CBK���#��{�L����SC0 ���:�� �&j�����|ylA���Iø�r��;�!u����]�����rF�+"��y�8�bi
��b��`RFM_;�d�?��ZL�Z,Jb�K=׹ꦢ����ҁ%`��xlD�̦4%�<�+>�u��)�~��X$�'�)p-V�Q�FU�qn#J:��>�3$�a8'���W*n$eQ�n}k�)�������uepvB#�`ɞ��.Q��Gx����|q-�("���`��މk�DE���8�U�롕I]jX��G�N�.1E����D�`28�����Lj=J����k'lq!*K�- !t�W���su��B ��_�;Z����H�G(=��/�;��2 �kf�Oh�[�ً�XP��ü�B��݀�kz�;j�z��}�+�b��w��|/����.<0�?c��W߮�ǜ�h�3��y_X�ͭ�K������.���cf ���"ѴuY�p�u�~>������d;�y�}��#��FJț�-�QPoMeih�!���c���f��3dnaM{T�ϲ��!_�<mq��{�\{�����m��;�l_�S=B��ོ��/=�>G ��k3�h
��
ֶ��U(>链PN����GY;�UA��|��*3(��Gc&No�-)j�&̢���1����[x�U���6[������0�ǋ|���r�Vn:;r2Z�V���@� 5qMd+�� �s����e��j����� 7����!�t�E�P%Թ���l<f�N4��3�/Ø��j�s�ۮ�<���C �p��%{��0q�;�G��QJt�Ԙ`��|��N��O,IyG�d�G����ej�0��d	��b���bw�	M�g����k{��m�E]s�[�����E��9��f� ���R���>c��@����.֣Z@%�6�G <��~*&�����1��#�և���"��m^��fl�������+I�*��VX|���+�$�ǠLGJu��10 ���w��, �V���1�Q;UD+f��\�G��N���D��۬{`ԩ^�,Y1�������7}�\�z���Ng�ʓ�����9�>[ ~n?,H�k�x?T����4F�z��Pc�0�
��?@ᔮc���!l� v��rK����l
f�,�L��,!_�QŃ'Л��l"�'$�$>(1�mqC3�} �b�h�1�Y�2��%��\[��U��w�,gr
#K�ޑW���!G.`���N��a��B�J� R ���FM�v��:����e�1΄����['��jI����rӢ㹷���!��4ԕ�lo4����O�W�e����ڬ�8���fR�9��ՈA2�S��_�p#�';��8I8Ďɜ���Z?k$%�>��Ŭ`	��-�q��m%���n�h�P?^b����Ww_%���*L����g�t�Zz���_k)<0�]ɝ��Ԫ����k� �-"r�yy������̟���<a��:�r
����%���|F��v�r`с��8E��:�q��;ۀR��W��]b,^��n;)ܓ�����wg�}������V4Y�τ�`�^tZ�	��/����7^�|l��*e���x������V���`�5�����%�#�2̏��R��$^�!W*�E���C�=d���i��D��9r]UdQ�	��O�#���L�QU1T�-�F�Z��vt�A��q�0����g�W��uL0�c�h䎸��'�(�3��ɠ��T���0��Yc2@�L���'Y��"�/|!�9��xC�c_2����Ո��ts*�\��ז׉NT]&��F�� 7�ۍ��j�xr�|���(���Au=_C&(7�!���d�h4r�Ҫ����d';�TQ�Ƣ�Hk�K�+R
[	B�W������Ϗ�W��񰜲�X�e1(^��k#�� b@�Jι3���P�A2}
��T��;KSJ��(�&
�Gw�Thv�iC��Ss+m�)	�W�t�^q�Y�|hr�2���d�j�ЎJc�{���)��:����$;(�V���T�����!�S �7�v�M}+��p�{��/UAZo1���=��Vj�gm��C��(|�x���:�k��N�@����6{۫��Se��M�������Q�DQe4�5��c9ƌ3����vRft �Fr���	�)�N��}�7����zU_X�҃uxb	�Sk,g)�ٹf�@H+����_>u����j���GN3y(��|Ռ��Xɦ��H(Cyζ�f���3�
�� o�y�n���H���j�XY�����ܶ��/JU4��=�} ���T��y�࠷
�Dxi�:x@���X=�*G����e?q2��;����y65�]�y��{�_:����s6k�f�T�����p,|Z�W|��oYϧOǜd�yaS-!���'��9���*(�Eԕ|�JOf��8�{w�]����3"H�n��p�M
Pƭ��J��t!�,�EAs�i�
�� �q��S�j���&�Xx�",��|�䙡OQ�Q��7��:��Q@��%哎�`��9���:�^��1��[��o��&��Ѽ� ���Yy�)��X���B4Ԏ��䰢�6�����%�q�X�$Օ�X��$�Q��"d6��c�6 h;�[ RLv ��{��զ���'�_4�t��������T���a��%D���a��r���<�������P�j����fض�DA<�(�O��QW�7E/|w�i �v��!�|=<^v��h�;��JG�����> bѿ����+�xa:{�;^�}^��(�?^�i�,�X�u�f��'&֞�GAf����C.�[+۴��Z���	#�Ke�VF��0He�$�x�GW��N3 ���/���c�$�n^�)�:'�C>�;�[w�	�d�[�����#���1�!{!]D�c�K�_���QޜO�ه�;{�I=_� C��%�X�@Q����A]U�|b��C�� ��'��Kk��2�Bi,1ݫ&^���=��o�ɨ��{u��EW�PW+��/���Ɗ���+sy���y���7|Ѯ�LN�"P��]�5$!@檗s��vx�8���W6����ș!�0ӟcf][���䤦�"�bl������d�#lI���1��&7�w>iU�����)B~T�n�Bj�?��}6еÛ#�������-Y�9�ͣ���W�ʮ^�(����M7��(A������ț_�)&yT��f�
��2��{��/*ˇ?wWh��#q�8FG�@�W�%Ԍ:/�
�lQM�<���d��NU(I0�t��P�٠�_�1���$�w=z����s�䕊�u���9�X��ad��V����3!�i3S����6S|�?�'�e��Z⬫ofE�Kh�ZyX;��l=	"����=�����uL���f���������������Rl�i��0���]���������	���Wɥ�4�������=�D��k�N�\�?P�r�>����V�mLJ ;߻�.�>���
�x������S�5�mĔCw9����AG����#�>&�(�8˵ǀ���R�P4���綂��lZq��P�y#a��/��6�;v3h�D�Ԍ�sӓӌ��Ziʞ��ۼۅ�$'�zc+%���S��׆2���Qt���]�SX��M�V3���m%�+P��2��d��X���m}�3�JmW1je=�6��}߷3Q��l�w NQVu��8&�P��+�d3;�tq)7�}��i�p8I�)�2�5�Ej=,t;��Wq�}����(����Z�tW�u��>@5T�q��$�Av]�9i�T�0~�hP���5U�?a1đ�RAG) ���Lt#?�.������6d�U�a|{N����/���,�ϜG^��0����!q =�ĕ���*��(�[U�L߭��A�[	�WMӶ'O��ݨ�}�y�H��Km�����.�*���t�Vp�&#��f��w�$<ޛc��YS��.rN���U��/��\���m���q�{ND�դz/�����l��z,����{~��z 23�cX �V[L���d�D�����){���H[?����y��'����/���*��`q<{4���΍ Z�5{L�;uç��O��-��(�ʳ�����Z�@D��DqsM���0&���$ŠQ/{�lz��!R�@�o�����:ZZ�X�)r��g\���D��̓��B ʢTp ��̲}�
x���*���-W�H��͟�	)-]���I������ȿ�t��Cۋ�rg�]
TaV&o�|�bҐ췧[���t��m�C�N*��n�i����0�#��D^b��f��3h�G.�G�����2�ϑ�1���Cx<m�6F�\g=o�箙���IB
����Հ��u6=�L�P5�]�Kރ^?�1�^1(6�.SN�����Mu�Z�9�k�ZG�R�~2��S���\���,Q�L;}zP7N������,����հ��L �,<�#_�%�$�'J(��i	��E	9�������͸*!S���z�	iU:���
�Y�
O� �c�[��7�L>��d�$��x��k��Y����W% ���@Ÿk�b�Kk���3-�d�yϷEg��J�"���e_
|�I��u[?��I�{�	����SW>��l��{^���%/�}�-'�����u�W�hw䐭BZ���"���O�'b�X��^����/sQ���f;��F���J$�QӗF�
qr��#��n��6n����o�������.� ��@�y�r�t^ҿF1�w��9�/��:k_�bN-�����Z@�X����RݡV�	[͠�[!(T���H�^]�Y��}�_�cd�y�p҂�������nA^墣
~ݔ����N�X�בZū�(�;�bH�L9�?��j�z�#����z���F(d=q^�}"
.��*���Ԏ_����"(�4^�6bhQ����h��������EQ�0�ؔ������@Y��|'����\��W��/F�7�n����]p�D�J<)|��ۮ,�i\L�~ �}�o�XEvF��#��Rr�ǀ#�£��J��n&� ڭ��31L̏.�����Tc���P��s?�!�����<��[�܉�R�w?��R*�0A΋����|�_:>lowa�G�$_����AѸ8�#�>@!L��<�N��aZ,?�����
ta������A-�S�16����'u�����P�e�n�}����~h��m���+�ǩ'6�8!<�����ǺM=��9b�}x~k�@5����u�hR�;p*KH��B\��%D7-s���x]x�y�+���,|9Dʮ��k�0;Y�rg��&��2G$F���.�����7%ܪ��,��*�}yx7��gP)�e��t�0�x݁E��Tc�p�
�H�=lB�R��������}\O����u_��T���%F�7 �#k79Β8��[���ѳo��f�$"��yl	��y6k?�����P9���6=�=7�Ka{��W6Pc�4�l�=~��D�C���m���e�G��h�|���T�c,����;ҳ���8���CZm濚I�	�ƪkу�������A9�U�����gK��IHםG8�]��(¡@F��'��u˻0}��s��r�n���ͩW���J�X��6���_/t+.����D���s��^�#A��\\�@:��:�e���0z+uӵI�y)�lO{�穬kڐ8�����gӡ���g��A>P�⯐�(J%�$���d��"����ؒ@q	�qĜ	~4��L�߼�y?n������0fK�a�;��['����Эi�*� �>�����Hsrn:m�Iಆ��&��TE�~*$9��3�$ ��~���[P��<�/{�I���І�rYP�7r�~t	���{Я6.�u��"�+l�ж@�m��[$(��E���P���I��ºSRs���=\�zw0�֛��ٻ�H��\M�*`&S8"2iժIVFΙq?�C������	��hCV��_����#�t�|�H'$���_�G��N�����,�@3x�T�����1]�Ҋx�H��Ɇ�3��Αn@ǌ���GS���,�:{N����.!Q�Ft�����?d�H)�^�L|���Y�h�u�/n�ѐ*�
�Z�vJ�g��º	�e�)u.�j&�;?{�N��ɐ�Jt�w� ��;4n�_T��X_��S� �D��L3N&�K��8��c�{����֘�Jn��0��C��ٓԖ���7E����� V ��������]�ĉ���]/��<R�KIn��kNR�y��+�\'H>�C�I�X�km{lY0��� #-��w]񗊏�Ɗ�~E��A�W���w#7�ZVAu�5_�>G ǰq[ȴh �K��v%f�Se�.��x*`��Y�6w�;U�br�9Q�S!�����?DcUS��L]�=��Q�m�})Y�W��^��
U�T���jϛ��;��SB���U z��8K�S��$#��g�>̌�Jə�QhR��L��N�<VԴjq%s������ ��>�dI1�&o�6v��c8����3�UpJ��5(m�����-�'^�52�`y�ԏ�������Q��x1��Ȭx�v(��K3Q�(tQ�ݥQ"��K��	M�D�4�9��P��	T�s�Nׁ_�Z��š�K 1wLtK#���v��"$f�q����������^ob���8b���yb��G�	����&�N�aA��
����[��ł[��2���A�h*V1�εi���[�ɫ=3���mBI2�I��Ehb�e6FVMV`���k$T��.Q"����g�'�,+ߋ��|llr��Uf�,���T�EG�jH�̋|�?�Ґ�6���x��7�n�C�i(n��¡(f�P��QG��ӾJq���d�=�;=�m�=xb�6��	O�i�������7� �Q����d#p��2��2�)xZҕ>����hJ�c�K�s~�e������5��C�{<"�����t����?��tM��P L'��z�zBy�����D�Yu�����b��V�0�Y.�)vJ�ż�m$%,U�L4�����%���6�<K�'��W���Q��x�~z(�O+ۤW��o���ʇ���x_�^����H��m��XQ��|[��:W�X��Ǟ��᭤)�B�Ғ���
OJW_�:)NXѣ�H��\�Q)Kb�}�ڳ����U�l��	�T)x7\e*Ic��f�Q=��)0FJ|�Py�u�����!����>KS���q��s��3��.l�}�״߽*�B��O|D`7/�j��:}^gm2�@ޟJ6���+-�����D�K�C�lx��܏�����n���\ׁ�p#�:��dk�h;��[���_J��;�)c�]/Hʡ�Q`�E֯x��rk�^�jT�A��j
9M��G��{�E8&�P���=[�C֦���CM�߄�_X��).����i S������o�l$`E�n/5Z����6��\���n��t�����D
f���v�'Α�1mZB��aA�=��v�
��P%�W#���0��E���+L���J�������Zn:y]>-�á6�=:�φ��ޢ�.�e4	��-�1�)~͌C�Y�҄�*Vq��\����D�{��RC�B���q|J�� C�'ȁ=^-p�n>�u���(c��B�Wb2)ߟWF|,��� Pоg��u5x�n_]
�EAByGH�V)
�����84r����1�q0��bƑ$V��^���L���E�.e�����&��G3��l�_��%'5B������7a�*1�:'���b�	�uN�H�������Ű�YeE�j�k����[~�%\p�������ox��$Olba˃_�'���Āk5n��	�YM	�����u�c5�A���8S��8j�W�������;�@}�򈬽')qkIkҖ�JvߴҚ��Xg�����r�drF�5�J�����Nա+���f���Ixq�,7��'`�e��h"Gn]h OkD_�˲��s �vp�W�?~S�^�g��BK�t���GHJ�;"Ɖ�@daQ�+�A���o������w�o$1K�*-��.?���֠H�GvNϛ퍗����|m6#�������W=Y���	�����!�v���j��Vj��&C����q��|G�λ��`5E_ه�~�$¿��t�"��S���޼3��yK�]��gDx�xI1�!=� ���a
\��ڴ�#�Ρ���'՟P{^w������~��Y����0����i��)>�Ur0?��_���Y��g��L�&���QӯW�'~�ݠЛ�Ls�R;�#z�&It��p`&hbve*p&�q�c�q"`�っ�U��E��"(G(�[{�@cg�BZ������b�A7-�+/oL*t�����D�ÐH+J͞Fy7y�%Gdb�J�㺩��4��6�0���Cl>(�0���'ū@B�F��ET\�q��[�	�����˿�Z[t���Q( 1ͱc�1��V�lՃ�˹��Nw
��Ts�q�gP�L�_��am��X3%4��<ZxoR9߅햼!�d�+��*t�hOHa���о���&����D�,�}��g 5��D)���6f�,�S�`��zcq��I ���}���k�Ԯ�Y%��(}ۋ
,kJ���X�pɿ ˊ9���i�~�:��a�0?w���CT����|�8�2,�yi�Ľ	[���(�fU{�Ip��r�TxMo�e Y,*A���N���EcW��4WA�¤J��*�-��>Ɯ17�w!G�W3	���������/���
F;T��f��
�l4y�u�Ea:^"����@��}��+ao����LP�!u5]�O>A��G,%�q$�
�J����c}\���f�ZY_����Kw��}j"WU
u�아E����q�8p���x�L���՛�W�9?(C�1��T����n�m�Az'�WK�o����s��R�m�V�q�\�΅���Rs9�"6�6��P/d<B2���j��I�W�EH�U��*�+v��Ll2�=˾��Ð�y^R�xЦ��$���hZ�_�𣇪��[�V�v�}�e1��z"!`�ʶ �:�2d��]��;�oZ�� r�~M��⒭.�Qj�!��]��S��=�5�E!}+���q�_z��r+��s���L�`�e�kg��Tu�^�o�-o���{�m��N�@D���l\	na��Y6�F�g0��0hyۏ�tW!��E^����H���mZ���'E�<��{:���°���;�!�������>`@2*7����j)�qԮiz�f�t��;��G.���d���6
4� ߔV�v(��XU������c��A�'�ٔ?7Q���a�S��b��_Sw5���fy#���J'"�r/�4�^tv�$~e3�#(@DM��l�Y�qlǈ�'$�e�(���7P�8K8ݗ�}b}$ŧ�%�7��"l\�� ݴ��;8�t$V�G}��!���;!���5��Z���H�) ga6~+�x�!��¶�J�A�3o��XV���zƎmxT�`�s��e4ڃ�r����ڮgXJeH9Ja#F��ɬ��#�����4F���'연��2�������z���ˍϨ��eɰ�L��w6)�,K%�����{�pdl#1��-.;�{ f��K�ڡ�ԱO*So��ˈ�ka��2W	�<��s�I�bA�>/3*Ѳu�<s�#Y��P*w%rR�oB�C��$އ�uoW`�>������(�$�5�7팀�Ԏ�"�w
U��Ͱl�D�e�{`�8%>�1,��ܙ+R�k��<P���{��̣��3��#/"���b��+{Q�͢^�	Ei�4����7e���lQEX%s��:*B��c{P����P�S����aO6z�?US?�ݓu\�7#~#�:9~n�F�/B���k\X��$��d��pS��d��ug�������M�q�ͩ�=F������?:)+�\}ӄlqU�<���j�%c�ުt}:�o�w=ߗ�W�!#N�?c��M�q����MY��@�D�|l3�8ɾ���t�ϒ��ҁ���� LK�
���뫈�
"�pt�����Z��r�l�S���~D��E���
��A�=�fe�1��W�]�5�n�	�|\�hhs:���n�(H���?T���#nf�+�R�|�]��]��hW2�K�{a��*E�2�&����b���1�Knv�6�ƈ��'��7�Zj�A ɳy�|=<�� %	�X+:���&t�����<� y��Aljy���DD�C�2���l�s%��f�a�H�Q�hn��G�eD��M�FJ1��Ƞ(�x=�X��C���eq���UxH�L���� m����N�a�q�����k7U��1qF���w����cw�m���>�6��Ѷ\�%V��U[��|�P�@�f���$�0ݽǩ��w��X_H'�Ђ�T�{/U�f"�8F������-��.O�.|�DK��,6B2��Qi�Z���|Q/�
i�]爐񶁾Z�{BC�Y�٣^^�
��$z8��o�wL9�$���10�ad�ra�~٫���	�ڗ�B[v���{�'�I&Ï�,��CΌ������>�C�Y.]�^�ӻmoZ��R�2%�}q-��'%n�c-q�C�ݡ�js��!h��)!-�K3aX�Ȏ���<n�L1V���S�ˀP4G�����ʉ\l~b��<��B��p����c9p� ��?I�v�����;yL�%��8ceL�!���߲E^�B�y����$K��3K
��(k�Eݕ��4�{U����❡ ��!�7���6�����)�	�7vbZ�ze����H��4�X݆Fxɽ��V����Ȉ�Eu��2R@��ob�n��o�?�h ��Ev<��W��X������w��v;��[o���3 �k [i�y`2��0�����*{s�	D��i���"<�ŠHu+?��M^������4��롓֩_H�v�jh�d?���`�[��L2���U��0�M�����.�῟S+*";�(r�����٩ǘ��"<���	�����&(���܈1x�g��.��B��@�!�[����땲��\Co�)�@�+jؖ�c��K��vW�9�gbB�'1ݝ
��(��u\)�x�1�.�_�%C�w���0����2���G�m{�g[�pi��>n�6�z�l��[7�<�@y�%�%�7/fI^7�;?�;��W���¹'J�R�����v�)�V �]�)F��f��i]�T?_�1IEYi�k�&'�m�oLغ7L�b<�##X� +63�������X��+5��n����2���4�4*t�M����G��TӘ�y'��.�j��&�i�l��Pr���6Z\�dR��jl�6�1�R:Ռ6�.�PB��A������9�
�O,���=���q�J_M�ȹ��9�����#��qٚ�\R���B!���%fɪW�u���,���PӪ��% "IA�՘�C5�d0S�S �m�	9`��4ĢuƊsFT��[�;��b�^袔�m���*v����t�Τ.����\���e��NՑ2o+�g�"�hZ�K]�^<Ta|��)�YC��G��R��3�?M�R��1p������)(s�8Vs�ܦ���?^0�r����l��S��d��c�e)+�(����� ���w��:��C��sS@,����>�T�>���P��_�������ےY��i�W$�?6K�)7���[7;�;x��m��Bŀ$��Q)�z��I�=���&�>��Ա��)4`M�cM~7�N �ڠ�7,87W@�~�n�#�]����=y��LN9���R��Q���
oL������_w�����W� 7���u�wܜ�9䁛L���H<��܋'0;��#b_>�����=w8���J�枾��˗Ϗ��D��o�'䃢�����:6�$�-=��q�����5�mr��-X������k�[8ep��e+3�u�"WK�m��A<�^(��d�enD!n4#_���j�t�o1 ��bgVEu��]o�+�\WV�>��� y�V�|f��PGGx�G#�^$J�s%�NZ��I)}/1�y���a5Z�`df��u�*
�$��=��:&����Q,�2W���)��5ǳ�.G�Y���#��r,6����]q�M�=4x��hr����q�l�r-��ܧ�o��mIMMu�ëp{!�&�MR
I�ۚ�e�̞n~���L����m6TEDz<�Yn��	�K�h�� e�q<?XI���HF�d��M�"�����<̖ۤ�-`��YF`b�� e��.����=�����(�����ѐ��{e<�0����E/h���2�J�8����x�$�f_���7o��e�s8��{��6�<�&�?�#odK�H�Aj�e96�G~߻�mH���%�>��k&���|0��������S)_��R��Bo	v6�+O�PV���,���l��V�[�ڭ�)%�Cɺ�S�Xym��됮bR�M�D�O��l���,R�H6!�ꪨGϫ֟��հ�8qdkW��UL̹�$*e�q����]�s`���f_�X�HZ7�@J��/	Ȅ��(qw��&�����Ă�tR��{;���cQVA�L��׌߇�����<��.(��Z�7Y�|�=�������^xLC{�)jc�N�+~��:��c|&�;փ.��gƮ���զXI��E�_vj*�-��V����p��O���δVw�M����MO���Z�v�[�Gc
4ķ�E����[���B0�Ǩ�4�*�Z���4�r�v�ޒ�"v�0 �4I�{s2΄�L<C�چ�^�Ͱb�qXw)��_
(=p�cR��#����o���w�)���،��f��l��[��4wp�s�J8b��h,�X}4q�oAh6��U������Z 9D���Y�����Y�,��U=bVd��SmMk�`�aE�Q N��̅_V�����k�WZ�Ai%���f�[8��_�=Ш!�9�_ ����5K=nީ�2S�����K�5p>�>f2�g�� @c
,]1��T��:������f9����8ܰ�S�eA>���BDϬ4��B<8�_I��Ob����C�6���z���`��\zws$!&�6�a(
��E��
���,x�j����cnm��|;'�A�s��M������G�7�T]-XyW	Y��`�c����)�Ϗ8c�Ƶ����O�D̑.{f7���ag-ﰛ��\���ag'�/�|�G7��u���p/e�m�F-Rd�jb��4X��۟и�=edO'�����Ω�7��7����撁3JW�M�O�R��p���R"
`F���Dr�f������>_�<G�m@��YˣQ1� C��«� M�<�����af|�c0��L����{6,�N`&%�"=Ixz�t|Z�A���A���h�Ő���� tu�
G�J���YkO��7����E/�r\�fƼ����
����ί ��~�O�G��Ƅ�qwP�P�n�m��-�����4���k�ʡ��e��_!�![m��:Or�9Ɛ4ݜQ7Z/�㠸7�9u1��M�*�}"\ eQ���ʜi���8��$)Qz�ژ� س���p��y�Ƥwn���m�*�=Ƶp�Х�/7�OP�?A$�R����H�z^����p�Wq�ph�;
�׺]pňM���a�ŢۼL/�	���e��p�n����Oh"�NZ�;ύa�+����3q9cי�G�*�����?����qO�PБXA�ٛ��pĀ
�`��\�L�#�b�� l_r����G'������#jj������g�C>}��^D�9�?���|���j{ �?4��(���m�=�¹��׵�%�پ9��d_wC �s�L6�_�B���w�ōz�r���Fa�;��奂���=�T�j�Ic�#�9���^�_��k�\�$4�3��*H�����rɛ���ߘ������U���%(�#��*�T�F��i�"ǘy���ج����q���%���p�Q㷲KIP`H� �4�����(��&���h��G�K�d?���(���
��}'[��p-�������o���uz�]�c�ɇN1S��ߴ���I� %GF�8J8�u