��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&|J� ��
�4�n�]E�V��۪��.]��z}o?�I��O��dĄ�*SU���A~�e_���x�tM��|��Q��g��т�IHo$!x��j&@���K�swU�9Ϯ����(L�'���A��f�z(�n�C�D~���@�'�.����bܾ�'��h.4��`Y\���;O��<��(���LM͙j.�':`Kěv��HhHn�OAD)�<���lP�7�-�z��b�ݨ����O�6D�L�e��Q�j��/�n��D,��c���W�`��}���O�PGh RB��,�q��z���*�>�o	�Y�c�Br����:Qڄ��䶧i���Е�[*��,WX���C��u��^�x��q�t��@E�E\�@n�{�V��'1�u~�Z[�EJ5!�1i_B�F��eBط�/�	��V���Bn�eAHC�C�����,��єM�q�� Oz(5�b���GHث��_��6��v�a?w̪��!OK������xյ=Z��MZR-�1�P<[(��^f�n�F"/T���uhPv�kl��Y�W��[6pC{%ak��_�4��el�:��F	��)]�N�Q�8n7�)s���b�Q�o�������K������ȧHKD����ʈp�=�ٽ����)�gdn�J���Fb�5=\~Rt���;e�ݸ��0_��d?��u�*UTi6�� ǋS�m$=·Y��}f���2�S�J���"i>��|o���	�6�S��=����/����|[x��l�,�ƃz|G	�Ҏ�Ѽ_2*,�̏`����k�=nb����Pu�{���<����������'��8���q��@qv�v�w	�4�?RO�m�cl^(�� ��S�Q����{M��G���*�z�۩��\�5��G�ɺ~��c�U�u������*r%7`�X�tiQ��G^�5q�V�u¡��C�����Q+�X#����Q����-�,pS��Dh��X.�R��\HshI��F)7ȉ�۟3�㒋P����f)#Q=�g��\��HDիZM�mg$@G�l�X��.�.�|oC�`7��/w�6���e���¾��cbd�EUd�
:�_������Q�~��%���%cPfI���~��T	��˟�^?&��q�̞������T�ֺ��.�Y��I��T�wR͝�(Ӱ��M%~4̸�t���y��v�U���I�'¸��Z��wY�Gr�>���*�Qp�P�3��{_l����u�}���7,�(��H�rP�9q�ϭ��-���d��s�����ܩ��(�Z{ɿr�X��s�j~As�TVXi_�������V��v�t*�T�	�� �CB�T7G�V���m�L$:_��Ji���)Q.g��%�
7n�F3���V��+����d�u��p9֍���Ł���q��D���Y�"���Q�2�W�p�Q�c�@�fe�S�䄋Ʌ�k�MZs;K��]M��[cU't�"���
?_B�_�!������5�bYH�%m��+��k�ý�����{����d��U�e6���B�;O�x�ET�F��+�L�����+%�W��hA��H,��ʗ���_�J>4� ��g�L�7$ˊ-c��=�'�ʰ�ˏEo��(�E���z���.:�T8��1v��>����n�$7�D��z�R��MDtN���phGE�r=i�F1�a9i��	2�wdtq����wv���AXe��G��N��5��>��B�\�P��o��;L�����<$k��ݍ��o�j�Җ���>�y
Z�f���5���\*�2��CI�/K-�"��g�W�?��ni�����~?i���rƵB"�Z���eX%�@,����)���
�lUs�(�&ث�k�`
I+U�^Z���D[�ם9�*��^�e#�#zB��[����VoA�Z�<r%
i\���N�Dhu�[`����(�;��m�%�+��E�j��E)
�*bU D���}� }�������N��8�f�8X���N	�M��j1
�r1����W���n�o��F=Her���BV���W��,C�ʖ�9��a��X�N��+@�x��`��B�wJ{��8G�c�u� j�I����]98��6���6���Ơڃ$���n�͚�t�9�<[0��r�\�K� h�b�ŝ��AI��;L	$h*?���"�����4져���� d�����R�blj�B�
�M3�c�5��޾\��� �ͦ����f�Tb���:�t�r*�#=N˥�����2���Ҳ�b��7F��p��?Sy5��������f�V~N����(ⱓ��gf���:��w�h.5�My�p�_��3�
����]�o. Ʒ�����><��d& �X�(W�Ւ�ƖWI�`7V[����"/�j���!���qŕ_!lQ���^�hꍭ����]�%�w��[ڂ��02B��YM��G8�Зʼr�x���	w�9��]b�|-6� ��R/S�A�t�L��BsyB�o!���H��FS���=g��ֿ�p\6�h�� ���8u<�)L~`Z�'�5����@Ņ�\X�v����G|���b#{�l�� ��z[(t((���AW)G4�bu��Du�N�\qW䏖��*��b���ݑd�x.�I�M�IB����ES>�}j1i��P�'��T፱�v��KQw5�
˹�m��DN;l����~��|oݾ1f��n`#m��9 ��`'A±G�U/$��Z���{�� ��W74��;��h�{�٦=�OТ���/��<�5���BU|��ً �w�h\}#K?��	���@� ���药�1��/뭕]�����fި�p��gF!P��3ּ�2��T�f�7��7����l�p'�y/�&/~��H�5��@i�`����Eߤ�o=Q���J#���.y�6�P1<�Q %#����Q�Vl��"�+=H��=��&�(�=*1�څ	&�=�P�-�4��l>ާ�V�L\����X���/4d��h���Y�� ��PL!��|��Ab4R�V��1�yX/Vtx;��^N���?NauC/zF��|+�ɾ���J�-r+��d>�P3 V˭1�r�+�;�k�[�L�1teyuh��m�}���=s�$�qv�\"Q��%߀0v�Q�7y�=H�`1�U��0g繇i�'��7�m�E,���R�G"e�{Iw��ziO��*�8��)��_YK����퀠�?:MMC��Y��s�wLkBWK>6EP����*�ɟ\�-��rc��k�׭���9N��
�9ף�x��ݛ\j �QV�.�N���f$~��:Z�`j�<�%��z�7~y��BN��Ģ`�w�6�FԽ����� �����X�\�_:)��"��<�0�M����A'�>g��-X�#���	�m�I<y$���N><���J"Z�<Q/I��^�K��{.�[��א.A"��c*g�/�� &��ts*��-d�)�C���iA���oR��Y_bi�!])8�=ĉ7/o����5�`��v�[@�������ܖO潀%A�ԓ������n������M�ζ�l�[�tEf�l?�D��4@ޡ�|4	�«FUz��z�~L8A��� �L� <��	�g	���/3��<��)�����m���[�<=i �مv�(��q;Y�-W�{�X�'�=
�õ�'�5$.�N�5���"�ٕV�M��^{#gf�5�*~�'�3�O� ��o�����\p$,���,�\����~� �3u���<.�aO#%��l�xa�0�߅��%�'��N���n���:CDX%��r�����s�a��M⫮A�7��e���no���G<@6j�oY�A{���5V3���'X.SؔN����ә�E9��q��ђ�y,�'�E粈J�6:@���Es;���Hg�f���X����Zv���0����
�8��"iz�����ŁA��+��7RsѤ�_1p�T*_/��1H���VM��W@��� `��_�G���Ã���_Q�4�m�,���Z��1��V�.*��.AAܾH�l���g�?P�E!�W���Ж�׳�K�0P�Z`������%�&��[���G�4��F����g�қ����U��~8U�(�L$���ǁ27J��)������T��aJ*�͆���9������V��=մ mĆ	�N��&�u@B�/�=���	CƂ���,����)?j�tu���͗����Q3�NO�:x���a��fL�'��/�qՅ��z%� GȄu���rf�_M2P�0h�5/^y��T}�٥D�@O�����YM��ES0��+�M:dD0�5K*p눂]yJ�ܤ:��%�Vt�Z������|Ѩ��YD�l�a�Ð�R���� ��yū���vt(�N�^�ku��ƀ߬�?	���]��W`N1	S���Pp���H�(T�Fa^)2Z�m�>��h�$y:j<e�*�B�������x϶�i�_�5oQ2uV��S]84 �&��[�2To���"ղ%�!b�N����>S��C��>|<��/����n4ڝ	;�c�5]-1�_��>Q-���2��)����L.��k��粳<��Q�y͗�Pr7v�`��W����[pb,ĉ>7�Sۛ�.����&�P,4��9Y9��밲�&�����rp�fn 8��[���+�� |-i���m���
�8�	(v�D&E�� y��h"A�e
��އ�;�2Χ��/�$w�v���4�~�T2���B�?!���Tf�������q �IU�5�hӛ?�om[W/�$����&i5�f�����e�ǿց�Z�³G+D�����un.A�Lk�ҞkR�WؒeB8�l�I�\�������3�$+a�hob�Ӈ�'0��rY����_7��q��NZ1��ٞAǯ�~�.HL 4t��z�W��/x�����򎣃����eM���8���l	�Vf���K�$z�R�	'��
b��ں�$�ـ�����|+{W� �3'�6�TO:���w�K�q����[э�����;|���5���R�A�,��T9ɞ���b��NĆ�vx7���%��y=����%�s�G"��l��d:T?_��`����������tQ;=�X���AF��)�4���5���6R�=�	���)��wz��7�ͅ��a[���1
ZOU-���$�x*Jtֵ {ѝ(��Qp�4Y��pK�؝�ۜ��2ꀟ�}ռ�y��o�Z~��tĮJn$U�����p�$�l,'r�p�?_�v*O)��!'M��f��qXTޙq8������M-�(�]��7�$��on��&+y������d~�v�i�*A�[nj�͊�O�7� �叟�Z�Ÿ-b����/�Z����i
t��"��b�u���V���è���R�pֵ/#J����q K"�^Ƃ�S*���%�� ��7�>�`�.`1��w��Q��P?�8�L縈�}�:B"����w�.���h:f���r7|�)�(;v���T�d�[l�m��%.F�]�s�-�|l��R���OqXe����~q��qb��Zu�|��w���;o4�R圁ߘ�Zۇ� �:QQ
�ml[�\�V�Zջ͆�m�qr�U��	�W��fJƏ�%�D�1���#
��q�0?e)�v��v���^��o����
b��"�!s���
J#�۳Y{��g�:̆j���#>5���2a?�����R �pz���>�˖���.W,���0?=�0�(L{�w�܈��bAFx"%�+pߣ�r��S�RB�PI�:��ˁ;��G�Y�'u��I�Y
�V��X���	|X���v���⩊���@N��+��K.~�����D�1����:=�����N_�~�����&��B�(RQ"�9Oe�|g�A�o�q��όM��l��8�_,3%ʣ�0�����Y2n!�_d	�	4j��:���Y�������6��[� ͣǠ���s}S3t4u��爅�zq߆w�.���)xAF:j�$��`،��e Zz6k��̓	����j���lJ����@��%m0��Q�b�n�x��s/m�m��C�۶�[�"p���X����w�~�h��(�/X��FA����L�j�MI�5}҅~�g�P5^"��»G�"��dӹ�X�Z���fJ3`(f�I��ݍ��O�Y���A
H�9B(�ŏ{��.���$����;.�����f�z�˱���^�O��Wf�D ���V������aH�3��9��s���^���;P�Z���$����ߧdGaY�g <��`��<Uu��˩�p�e�7��B�4�,������%�2U�{�]^�^��8 �X8�F1���cl=��XS�GV����^�����#�n�%��2�3h �Ɇ�+�����0�:�cw>^�{���d@2�H<. �Y�9�����[W���O{���?)X[�ҮqCϹ�t@������ ���"˨��%:S�08�-�
G~��O�!�U�j@���%\;�hd�(��8�g�5���k^-������LN�^�Z<��y�w����U��[����Z#�_���P���_�v�X錭���~�n�g�����g^_*�%(*̬���>hp��g�`�+�c���N���N,w�bM�{�|����d�-�>L"�v�/�|:7%�߭}&�+:��
�j�i'�N&��G!m����K�$�Ǘ	s2RG�"�6���,��m��t��<����w!��2�u�7[��7���p�,#���:P�
0xK����2�<�$��Ё"����M��+��rp��U󣹍\6��V�U<�'�@�I��qsy����	�dk�Ŧ���K�q�بm�z$P�`$��k{�i�Av#��Ke���!3}&��}��Fs�H��~r;������/uą{�̆��<g��5�c;0�\��7�:۳BZ3�d���1�4O�߷+��8�zOn�5J
��`xD��5�V9^@3��	9I��nTI����R��V��S�Jcbˋ8@[`�\-���������k�鰣�N�8�m�S0]��>�a�{?���F�a��rA�����z��������� Ҋ�D�TV�m��=G�z[	H�~�y|����z��F�4�V؆�F1��ա?�$F�_��쪃�L�<Z\Tw��o!;��J\[��i�!K�2=p�d
z�>T\޺+STFl$e��
L��ܰ�d$��-��`Pupc�r��!B��\�YD���_�c2^�3�#���`�<ց/(
&�8���K]E1ja�No�7t�÷;YA�Fv��6�������f������K.?�u�5�h�H���F���S0��ub�uc�dɯ�l'�k8����,��s�G��!G�� r��Љ��B�1z�f�揙�f~��ܑ��6L;M�N� I�=l��`������ ��7��5d(N���O	!���!g�ׇȏ�X�_���C�"8^)�Xמ���0��0��;Sy��(AQ����J�g��6{7�!4Yϭ���[��� ~ >aV�����I�`��>�����U����ի3��� /E�/JC��c���f��Y�||��t�a�#[[���3��Zk|��l�H`�meQ��m���4�JU|���F\�0���vC^����1{E6���[%��t�F���������� �=U!�UP�p/֑b=Ӄ����ąJ�!wS%��jM��~���k3��+n#9n��Ͽ�"��x��g����ad�cz.��:����3�%!	���������J���-�8��Ѣ)���d ��
T_�p��hj�"khv�E��bkRR��R�;K��vG��)��$�0��;R�"d���R��S��ܩƍ$��xu���Ek�jK84�JM�v�w�1D�����V~�q�������?�*Q�D�x-A`�e�ЫO�`a�)��%�8H����A���������|�����B���d�_���'�����-#��ra��;#.�O��!� P{9y�؅�r���;����ޟX�[�5	��z,zq����[QP�hc�a�|�_cjhՖM�58�p�g���a�C�K�s��)���u�´� /�_�k��k?��P:�I�]u�"Jk���*������e3�5<7&2����V$�o�2�=���5J��[w!���Z��(�{��Fv�H�9��˦�'�u�������b��v���o�b����� �U�!����X�z��Z����2p���L��}���yނ$�g��j�ǂ|EO(�f�=���w)��Ye3�].�u_�(L�dT�*P���6�h�C0���:NB��B������r� "N�@�z�|�u0.�o�e�b򉘹AC�"���|W~���.M��"���͠����ulKř�� �'=��UF�5:���_����
o������|LY� ���Oh~
J����q��3�*��)�b��d�p5@��H##6�e���)��ٍ�_���G�wS��Qq�����xSliP��q9�G*��H}]�� 3j�څ�g͌����E��r����h>�G��"��K_iH[�w�[.ۂ�%捻$'��.��7eq촢��LB�\�c/(.�������?AHW�FH����ED3E����~A����ԿةE�XAF�A7��z7-KG�`����d�.�X�\H�w�Ц{�ґ̈́����@�uM~0:F�ݦ��aHM�=�	7!��$��t%�5�.(�3��j`��x�r
��(�t��8�~5{?h���
�h�d�����?�r�v�c���V\�-���M8N�$�*�q��;��Kq�퇳-��!ɏ8�̱*�����z�MD���}e��}˪=?~)���E��W,t^Q����u˃YY�т�:X��?"�Ŕb�}R���b�,��NnOܺ�2������Y����ؑµ����i�F��Rg�q��D���%�'s����Ѽ	=U�)�S\��$ꖀ���5B��G0B�� �Jd��s?⋂��- ������gD�}�e1�6�O��7��gQ#�̽�k a�?JGLn��}��eK?���� ��}�6��|�5��һ���f�㡏]�O��)d����T����hX�Ү+<Z���cN����0�� �"������+�Fb�:u\�'�a'�k��uy0��5O� �ɚO�\t�jRd����b��EO�Yn�A�I�P�h���ljA.2Q�h���y�iK���o(I0;��9���#�]�.���㝉��c�:9�]�.EH�,�D�-M�o!��p��'��~�채%=y��U9��mt W�Z�j��?�84��d��)�� I�Qֵ�ыA�%���RɲjÛY�غ`k�E���<~Dt�ȣհ	?�`֏X�A�t
Л�A���Ց��P�SX_��6�;gl�qO,�@�h��\�-n�<]_drk�GL�h#�9���nRZN���Y�[���<"�ȏ�HNq���BQkV�Lh���6����փ9E��q��|iy..pU^W�K=㦻�I^�������ꪎ������)h��l���d���w4�Y�M�H0�"S;�>5sA��8����LN�ରF~o-=���Ա�P-�m<��P�"���t���s��]4�/3ԚO+щUY�s�S�Ѻ�K 8��Q�ˣA^o�MQ"��檃86��_��B|+-
�~)U�U�uyTl{��8ΐ��&o����%���p��0�[q���=5
����H���N�hfP�LPq��D'UƊ��#ȥ�k�����J*~�8틗Rw��p�W�ׇ�����m�cUUS�D5�)�f'�g��_l?�\�Z�I�<"��W�����M����7�3O��7��""&�@r_;f^ৗf�����i�M~h�w�W��r�D.o�ٿȗ�t�p1��Xy�����K�{fM!�����i�0y�.XhTJ?�o"#$<�Y9Ef��!$��h�Վ|OY��Qa��q�E+�d�醗�LH��Q"��1��Xt%�b����ՖUC3C�7��ZB��0{�|w��C�WX�`�m$�C�S��Q���'�P��U�v�A[�$�Y��Y��7i,w^�kW٢S"Ũ�Rv��IY�K�K%�����}-T���b]�ݒ2W��A�"t��0T|,���E���RջXu#a�M*TJ,�^�;���i)`�,�y��:y���+Ϋ޼6lS
�k[�ܖ>T#��p�+N�g~$�,��c�/�'���3r=3Xxx���a�ɺ�9}R��h\I��K�ǉRP��(� uŶ']�JSН���]Nn*ɗ�����&��z���x��_��A�gq85�3Em-����Z�<����ʏed�1~U�����a=QU__��.�ΰ�J��fQ)�2�̉F��Xw���ĈF�Z�U�}�#E�.��A����H:��i���}T��/��-#��{I����l�A��H�$x$a؆Ó5����)
�@q1�6�.���(1*�-�,DB�5_����u��i?��q5�ޡ�dةL�I͙�p�� |톅��v$�9��~�G)��oo����B�R#�:�آ�[ib[��r��Wڲ�V�- ��:CӿP���hA��ϣwV�^R��G�)�b��~|]�M�8E���(��V%y���z:J5A�T��0M7t9��q�������n?�.AY������aד�T4zq@>���ÿǺ-󀟹>z���n�r� ���(���`��u�іQ�%\�X�s�Izu�������Zp��^.=F�f2K7�H��5�~����i��M�ma�4(��N��+*w����Eh�h�1�XC��%mޅ��B����K�&��N1��q������ �3j����6�E�w�dhi�Rw V��o
ͷš���Nm\��Z�͐"�����o�X( �߸!�&�M��^�4�$l�R��3'�R@�,Bu.46ݞ�^��f.��].�6����D�o1w'k��/
�?�Ӵ�3�ҿ�:���5[�՚}�`}�Wb7{�v��鞏,)�ؑ>8�YvM`��3ⰽ5B� y�����	(����.��B�
�d�&�߿�b�U^0�O���U�o?`�賓���{f.�<_3������F)��Y
��R�i�Z��-R�[�e~S>|���_��;[?ʦ}J���u�9�I.$p�OK��ͦ�,+.�r���7�FNY�RK�)Lo�VZ�~$�Q>�7~�����m����W����~D��ō���.���o˘�)�ȩ.-�9�;�ў �M��e���(����e��[����m>P�Z��'�cd�qk~xܥĳ5�B^���"+�h|Б�y�h\7ދ��N7T�v����w�j����l���h�����S!��Cȥb�?�C������c�(�0\H�7���f�$�0ìPva�U�������7 t���� Q>���&�
=�]J|ɤ1�g'	��%��D�<���ƮT�t��s��$�&J
�u����`����왐�=�1��1ih�vi: ���6yʣ�ŎCq�<�CX��(*��fhe�&�Ղ*��~�*�;�A�HU����+j�3m?���~��t��%�5|�����9�5H�j�[��m�����l��~�,嶔�8#{���Lq�fЕ��������!�fi��{⟷�&�;@4N��  ���|��PP�_K��X�Y������B�a��b�75�7��J��q�<��&�|�y�����l������w����Ʊ�SOS��Ї�c��]���4��\	0t�L��M���z��� MJ��$|s��i�?#!6}A�c�Pb�J��5�Pto5Y[�wQ����(��
u4�L��P�/��Q韷��(ƹ=-�<���N��J	 �����pd�>(��Ϲ9rhϥ�����A�t,�����nb*x���Z�v�$��ʷzҨ�뵑�W�G����h{��KS ������AE"F�ג����/�����F��j�y.���C�Wzp�#A+�*��%�f���U�>��p,O���(o��e�<�[��8[����mw$�H��dq��:��ӹlj?�(�y�Q�z���� �3�f���C��e`J�E�D(g��I6`���#�ndw�Ix�ś�vBF*9�/�g�W�����x-(��p�̯
,�0�^��Km���h�W�����t�M��Aa襜4s=��&���4)�_T��K�
��Úo^���<�Qo��7٬�g���C������A�QZ�U��a����Q�O�J&2�Ͽ��k���������"H�� ����������=����}g��Ӛwm8��K���2!�o�۸�J������+g�6�^�����i��L�S��iؒvNٿ
����x�Y�斕S��?������q/D��҉˩�0e�2�����;=3��΢�pS��R]qd1R�p[hZ�D��YfO}�#nUX����F���TZ�'�s��:]����ԭ�to��٠�g��5r�a��'<5���S^[;L�QP����UG���V�P?���Bq�6�j���g�a�`����2�o.����Bav��6�x�i+��nT�'�2a�W`�p�g��6)�4��\�G֑Uy`�q!ɿ�	~8}��][�8�]�.�q8��IT�3�qD�g����;l��4�j׳��n�A�m��볤�YZ�I�m�����:�2�+�?�vJf��
$y�n$�P�h̿i���o-�����¤�0�B��l�s��#q�eߓ(-2�_y��'��qrĝI��^סyB�F�m,[Aw�� k�8��,F@�Q=�M^r�/᪝��T�Vf��:7���o��)��Vg.2��L<Z�3�&^Y���x �z�ٝ�s�����bk�:E��]0�x��zl(��)���2F�+8��������4U�H��5wz�̲�B��c\C��񴓗;v����$��kH���sD�?^W�}]l��.����6��W@��-']	���g�Ħ�	`m?�0�s�:(��#���da�V�	��4��T�"�4�����~��5]� �a�"��<W�����MK�� ��Lm^҅�"�@LT����?*:Ņ1<-伏�\��CQF���rX�>M�w2ǜ ��94�����q��.�7�i����A�����Bأ�i�Xt&9x���!r��¢s�!�ʈ��,�
�	 �� l��e���y�����5�� ��N�Ӝ��):�Nv�z�.~9:N�����ù��)�1A�=��q!�&��a��5P��{�^�Xŏ�U���0@Ц�g��F�x���u5S��!�C��e����V&6��Hd����GW������NG�!N�4�OZ�ċ��P���؀B5���O���Lci|�~�mՊ���g.yq$P�]SǴ�8uN��F�(��$O����1D��Gb��}ԟ�f"�e~:��t�S\y��b �y�E���Ϟ�Q��Y���>t��zb���rm��V!��"��M�����Bp��s�������Y[�$l��8���-��2��d|��`B�ē�=R��$J�8���d�S��<�83�K��P�+�9M-lC�A���E]&��<��)I��m�Mo�_�G�0.Z6��dĪ�y�������>4ȍ?;�Xh���Q1m�Nv@^�w���ҷ��;��q����5�;��� ���L�X��� 2\;ٻBYmB��� ��H^	/>�j�A5����p�|�q��p,�fZl�$��.+���":����8�5A��Z��{Zh��gY��Z=F�z��Fv�����f6#B���%0����ь�Y<��{"���Ⱦ:��Q�26���p?i�v-HAT���/:m��Ż`���n�S��d9��v�^O�1��.��QO�;����疫Ou�ޛ��=��~���z݊��j7�rt1�ۛz���Bۨbx��Nŕ(�)�0?�0Zn�-,
�D>�,���?`t�=�}�[K�L������N�� <gQB���Z2�t�F�]�Q /�_73Ԃ$X��j�4xlj��,yw������$۠�|��k+k6v�ދ���:U|�o!]߄)t�7m�b��鈓��sp�gz0�Ct��T*!r��ϚeP�g���7T�L5�S �;E�"���Ġ�L�K�O}�"�U
1��ׄ������"��
3����������gt�]�������*3D�2>�sp�9r��;"6:��vUiÔ�������rކy������:�g����bC@�:8g��sE߽��@&����`p�1AHlE�q� ��$�&��@#��co�)�Lj�HP�H.6GX	�2�+A��aF(�3ܼ�식�4�*׭�Qu��X�U!Mx��\�\�Q�}]��� �um�Yg_m�q�ž�5�����-4g(i[}޽�|���#��|%�@
��i�2�^)���̓vx')C?'���d��C��7I3#�9�_�Ke#�0�v�[=�%K�zW[~ct�b�B�յ=e>���(\�e:ҥ�j��������Â9�q�d�8���ą���2L�����B {8]Z<quu�5�fqZ�HX	Ӳ��U���M,�[�s�+�-[Y�
�`dkn�p�r�ŏE;�S��5j{'鷃�)�(TH��ɋ&��^x3�� ^�^�E�t^�&/�SI����\���f��pj>���QG�f���&R�q8�*�եw�cEK�s�p���Q����_6�c)�G�G�� 6���^]�6�sU��h)p��<;1��R�v�p#��snތE�|���G�l7���W�97�7d+u��m�~I��^�D��G^ߴ�W����P�/
�T��t���<f��l�b�vlңY]��׺t�u� gJ�,9���S��8�|�5�l^�e�>ڊE?�C�Wa_1�5&��sKJqVW�	(-Ŏ�1��np�"�Ř@�����b�3�#�:���9����
��=��a��M�7�U�W����WlE��zj:�f����z�~����w���+��,,�^Sq=Xu�I#n;VzKh�o���1L���;-�8��f\4�cӽ膸�#���<s�G�Ԣn��&jm$���P5��~2��y��*ݢ�Tԍ|�m�Q��4��ҡ_B�-Mv@���\�(pY�صK7�1�j�_���?=y�`��VZ�-VɎ0![.w���ɜ�C7j�\J��s}腓���e����yo6?��,��Wq��/�:�qa{_���b�&?Ē�v�첞;���w+C�xX���T�<��Sw��+���V+�],vgą�R�#ՖgeOj"�����/.�o%�
O�E�+w%3�<s��1o�j&z�Mn�&]�/��L��[�q{��wTqZ�@x�\o�K����+�RA�q�݆���L�f[�T��-���w��7�UZ��g��`���'�x���:�e�IA�j��L���w�H���� x���'Wu���Meb�1#Ri/?-iUTT'�pX,�y3�:kk{�/�k�ꎞ�
 Jp�8�ka�؉���q��}�m/,�F�l�G!X!�b��2]h����'/S��|[Ѱ�h�T�H�?�i�õ��g;�IFr���F������l0��C�����1�OJ:rȕ�.�}��]I�nz�pP��!�x1[�R���&����d�|RP;S����(0��P���``Q'���F��	
����I��Y�=�WJ�ʆ�Ce�Cx�Pw	�U����tZ�Y
����%����"��d�0�~������>������l����XX-И������C�W�E�6;���$=<���ÿ�8CZ|E��n� t�7P���Y:@�_{"��M^��Y��ί)a����7]�U^q*�*�Y��v[�ˉas������~W��Ȕ�^u>n�9���4��wI�4W�j|а�o�"0�V��}<����"���jj���@����R �Zϩ�;���&ܕ�*�y�����Z< ����������#	��"��dOLvv	q�׽�\M��lϞ�Ȼ�rE�j�i��T$�Б�����m�S�*��*�����!��|�!���l�f�PK�d%#ރ;�W=��r����Ϟ��-��L�$���7z� �]֚����0�`��<Ȣ�b�ֱ�����U�4٦��!��kSA�e!�w�oxЁ�{԰�H���
X������RS�+/9G�B'�6��	�e�o�'��� �ǿa�g�V����!f�����Y�A����g!��.|�{��V>!R[���ݚ�mS��b﮹.��&��fE�!sTHEz�E4Rsqw��q*�b�/��ι��� �&��F���S�Y:L�JZJ�!b�Y��U��뛪'���:=)�ұ�*�����l�?2G������2y U5�73�s	�:�����>���4�,�����nĘ˝%���tV`�~B�v�?��/(S`?1a�\�S�H�N�@�__P�>��A}dx�!�Y�F{ʏ�)��l}����k+�6�܊���G�

+Y�=q��SР�9�th�	��C��:Uo�%�X�2/_���p�HqB�z���M�Z����a/��i��
���1
.ؑ���x@�CHq�X�,ޠ>n��oĂxT̜�,����]	T�*�D>��d�*>su�Y�%%d��B}�[�F��5#:(�F�ݘK�0Ѧ����p�X�lEF�,�/��✸j����z�YEֳCb�8K���!��"?"* z.!'�!$;�w]EoU$;ɲ_�`NR���7��鳠%W҄7$���0���rH[̒ɘ��E �_��cT.����1ڕ.)B�����Б�̒�[q|��5)k8"ܮ���?�{�í���6�Y���MY��>�$	wT_�4� w�>I{x�ޥ���QՊ�Hd����iā��1;���D:ɭ����o�R&�ĉh=Y��xG�#�h�3��f��s���W�"�@ե��d��Tp~,�٭�֥�v��3%�^�P������Ə��eǬ�1��Y/X�R7cC::�r��)��/#!Yp6����7��[��s~n'�OH��_KB�;ܲOx�4(Q]��>\�A�I��5�ЮK:�a;�gď��cA�w�N���A�E�o�����d����O�x9���n�h ����4��U�Ɠ�� �A$�^�(s2�2oR���0rb��r��UEm�_�t9TmM�P��e��w�+���*u��XA��m�n�6�7ܦ�h�U�"j��	���ٔWYXvV=�G ��P@������q��5�80�>�!�<s6h���W' �D
�L�<�6W!y�2*fP&��Ul�&՝�N��&����B�n�%�+)~��$��Ae�-��^�6�!~Ag���F��r��:RJ=:T�F���ؤa���[_,qM-�chy9���cu��k�K�5̐[�Yq5�5�jg�6P ��"�D��c��be���V�G6������%+�u%㟺]�OhJ,�����G��ı��<(c��b&I�Q�_ݵu�l}�/,T��_�J�	j���[ՆW��+�r#�X�[�u��Q��9KD�뼚r�E�=��q�0������Ȩ��M�����
ha+�>j�!�cr�5zL�Q ��p4qN� �0�5�� ��ʂ�8���9`E
.�,��G��\�7P(�S �4�'fbʸ%�^�k��<D�V�@u��U�d�����A:�������S�QH��`T���ǒ�����Ϟ;���1�2Ѡ?��R#E}�J���}mY�mAt��Z�O����9�+&>
���X	�uĄ��2���ޣD����Y?`��Y}��)KJ�_ʷ�R��]�F�w?��Z��,0>3}��h��q����R�{H<KN����a�$����i�F���4�b��SȽt
��b�jg�~zx2�����4*���k��'Y�Z��D,�rw^���E�L�z��&(,� �O3���E*�mrS{Dl	�4.:2�:B�9[�����O�)4$7K������^��jȓC�f����4�Wc�k��J=����c� �p^��zT���Y��Y��āܕ�� ����͚�_����}���T���hTi��6�6�����.y&�X�a�O��Ks���w%�p�8�m?��.��P�Bk��X�z����O,�`�|��_�K\9��f��u�D4JN�E�R�^u�)���P��$�q�$=��P��O���C���	�?~l]����3�� O�����́���}���%W�4�z�&ZH��p%�]�e�^�/�����!���]� ����_���V��c��?�A/?oʙ�4zui$�st�ڙ���1f��\S ��'5�}ԍF	0a6�萕�7��X�y�9K�� ��]l
��I>B8K��]�>l\�h�����۬�Ѕ��/s�c�8����Pc��y�[XZ�m:JV��%��$
�\� n�쮿[�{5�I�r�*����� �"�����rȻ��sk(�M�����.*��
�k���g�
^r<[��l�až�&0�*t�+^;�Ϡ�C(Wj7�ϒ�a��L��"A`<��M\�YCA�%
��`C�α�~��`C��5N��I�ꏥ�g���c@�(ʸB��ܘ�TX�ik��U�/��|�KC*j���+�/8�D���p�$'�kPU�{�u]:��X����M1��t=��~d<��T�VG����$���J�krf�W��(%t��\g(w~���>ۢ�ʝ����Iy�削R�q����B؊՚Zq:o�2vJ�^�͖��2�Y�^	{U��@nfo�џ�������_�>B�N�60�<IͰ�N�� V+;�*h!ҍ�c�,��`3�s��e�;6����׷}A�" <k:ˏ���Ö�w���fB�猪��)�Fy�|���ë
i	��P�e?�e|v�w$����� �����g�}	��1Y���1�
S��2'E�a�@�x2�yXFd�L׉z�1�&Ǩ`��uC����X��d��8{κ��su����5;4o�ۛ�4�{{�(S�E$wʣ��+~[��c���d���.��B�3����c���zW�n�o���*�7���*;����k�(�E{�f��	$��9Ce�t_��C�s|W����8�$T`�����R@ �	�����Dx�R�`�� �<��!Ӷy���,���^��Y@�����Ӓ�9�T���2�J����=�����^�5a�5bͶǭCt����
U��&��>c)�}燝����/�rꠗ���F�B!�1M���Ղ;�)��;;8���*_aj�`]�&���q���Ffŗy�=qx�j��O@�R/���"�3��σ,x�&�o]����b��31�d8M�.l�6�!�a�5��r)r�n#0�_�?F\ɒI9�(R��"!�_ٹ��� ���F^�v,H���l�&nji6�Qu#�d�2�����H�-O"�c�8�=a�ц)�:ӁO��u@$����[H�#@������ci{���(��9��b�F˻Y�T����^�oV�|�n��.�D����C[�ݞΚ�夎����'660f5I�Wg�A�΀���ڙ8��y�@@9�o��ٴ�K�p�aV� ��>4������<��|�g��8��<J�%nj\d���s�J?.��1���>�!c�K�|�{�D����e��ww:k��r��/@����A ;K��g4��GX�t�N��0h��	�
>���y�ЊV�g�\U�CW8�����-�sCv�bϧ�J �h���S���g����ʎ݂g��R(��j+U�Kn�:��ʞ9Hܕ�����KYꘟ3�uz2��|M�,Lvc���Z��UNI��w+�@}/�fU�<�5fN���'��;;�Q��1e`���+3���5�N3��3k�#.l�aL0b� Z6�r�h\�|���OE�`�I͗ن'�i�uL*�|�<|0�zx����S�U�s��]������#����>���cnMVH��OEo#�>�;˰��]"��bk��D^��U��}�B�Up�U�K��xz*k�F�6�B�]�9�ڤ
�Bme�/�������A��̷=���
p�a�� u�s!���Z�J���N����֘�nk��ͯ��Ha��u�������x�t���~zJj������U�aˌ����l�j�il(����k�Q�Y��껩��̡/����9����J�Ұ�yC]�C�����ԇν='4T�C��ud��9/�q�]�=2�F7;�, '���2���zD,���	����䗯vU�Ds�XR��Cw�����g��4oƨɌ_�xi�ct8�PU�l.B�{B�6��X��b�C�4M-0����l��wQ��j�ҍ�L&l���j��1*Z�;�8U��C���/�g8�vW��v;��Ϩ�����w�5	u�߲�~�P��*fc��\�}<r�ֈ��U�2sB��]�Z��/�؊�3��$��i^�$!�X
���Z���u��OL����0f��CɅ+Ӂ.��qJV�jX�0�Ǯ�ĢB_?~#[]7���#�R�I3�A���C�����U����=���*�&�#����9��T#�$��L� ���v��&��vY~�d��t&��Z�B�;ۅ5��R���v���Dj���{r�Z�ɿ��W������/B�w%�&G	$��0�����ˡ	�텃h�6^�o���'h:YDo"ͥ5]��g1��7-$P|7���Y��?܀�0L!�5W;�Ŀ���W�[�)XC���+��_/Tr��3+���c70ө�˼���QָK�PN��n����GU�鷃�� ���o�Y��B^@]ݙ^���J���'<���c����9��o&ȷ��h&�����(�W�#da�jA�����h�B�@ÿeLH����{ϔieӈ� 5d��$eay����_b���K0$��>u�e�����п�t�.-���*����f�I�	u$ț��m�A���]�R���pL��FN��(�؇M�"ҥa�H6�CD8�Z��P9�e��5�f%�ƂE��n5���qn��~�^6���T�Uo*Zi�`�/J@���ո���p��E������dg�T�WA�]��-��Hբ��A��~_���}���7�(��d��J�t0��h�t���c�7Iվ8�����,�:Z(�h7Q���$�g��U"��~�|N%�S�n���C��O
�?�.eY������]�w:�o��� �(o�H,�rx#�B@�_\ΰ�����y㋯��?\�����<��*����;peK0W>��)}��_�3��HWH�"��x��*"� �#��^��z�-F�R��Y�zʂn��g�ǥ}Mce�J�Co	6�#�ӐD�Ł�"/8�����$QPq�:�5UR�����M6s&�{���Ƽ$JjzUl�^xn��7��3�f�EI��[Zb�qa��w#�$���x���g��Ub�G�w-�����w���`���!$�z��Ǭ��a�Z���U�[{VֻZ5��f�é��7���GѢ+@| �������la�kэQh{Zzt|��M�<���8��?_�JDU��
{���r�[�����4��E�Ö�����Bu�b�ɹ��0C\��r�{�" b�"�>�$�7��W�`;�լ_ų���;��n	������,d;B>�18��q_a�\9]�n�H�Ő�uT�:��8��޸��ə�8����0�����Qj��i*4bc��l��L��ޱW�2���׉WQ��i�tP7'�T�J�s�Ұ��l��i���k/�\� �M�Í8-�;T]��e��U����w��8t�2	��]+��|�`'���c�6_S2�5a�?�]Fi��`�u4��H�S���6���g-��eZ�E��Z