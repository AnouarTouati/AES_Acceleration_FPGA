��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���ohB��爾f�HG�g�,ג��XD�_I�v��t�n'T�j�^��}� �<���[b��Ą���e���*�9�sV���g7��R�T���m�F�@7C0��Cb�, K���$���U�ŁU^�*�ƤlKC��inJ|�e�-���]g�~'��peG[_��c�97�A$�u��I�_ػ�sؐ�Ժ �j�]�G{�QJ�`[!�e�TX5`n��'�H�`�b,���${����$1y���T/��ɭ��]"h��/Ȳ{�����:c�F ᵬ��o@X��3�)�����,�#��+7����0\�	a m�#���N��ZN,��3z���xa܆_�ĉt f&�{~C�����b�^��oXZz&�|$�~�)X��$6	�w��V��.�^U�&͊�h:P)��R,à�*L�a����%-H.��$�?A�Ӱw;�-v�7,|�N"�l{2t!�o�Sk`����@qC�|�$e�q����"�sB]���樻�߁Tm⩡�
%E�mLd����I�.����>v�ecv��X���z����:����Cx�=uw����H83.D�o�w���-E#G}[�u}��+ O3]_R����4���p��O�w�dK�os��j�H�|PÌƩC��E��RB(I�*�q���!�I�X�(3n��U����{�Z-�=A�F{s�aJȘ� ���]���qck��~���w��Bs8��;�j-NзJ7:�y9C˱�{>��ek�D�gw���g���� r[QGGH60p�n�J��k|��܏��G�t�D^Pn����O9��d��rU�*��*6�Y��{s�>�mp9�~
 ������ꠗ7E�K�3����1��V��k��)gk�X��i��vx�@�qo��>���o���Co�R{��V�{ep�֦��!<>�[0�
}�r��&"�d�D�% �uv�}'sx�#�V��{�� lFd��H0J~�M�C%U�J��'�Q�)�ġ��`��c�<X>R��>Z[�����<h-���tՋw6j�	�yJ�9�z���ӻ沬��$�����>���fZ�F5�+���a�`���O͑+��
c����iHԽ��HgG-�Kx�m�1v���
#��.=�
Z�qS�7N�5���1�ϑ�o���J�&<P���=1M:��>� �p�Z�
1mB����5��X��,��i�3�0�fȞ�!�Ԟ�X�����'��qG�c�f_�h)l�cK�һ�i���7L��ƛ���}	�E��	�(������o��t0	q��K���W=ub�y�v�����f�񘈕Wڧ=�5+�c�λ����%�g�����F�X,� YX�=<���eǲ�=Z�j�pW���}sJ[Dhl�y�x��BLM1)���/lXT���Rn�-R[rQQ��`P��P��ߏpU�����ɂ���|!�>�^?�}A74��	�7C,};���|1�` ���S��K�;�گ�S���yȈ�-��+�����}��&�J��*�o�Rϫ1�j���.=�T.vK�&}�.�?o@�'����ƭp�]�R�+�=����;�3# \}�)�f��*� P�7����|�&���s>Z���]y�;�ò��������P-y�M����[�D��W_�c�3]�ۇ7��I��ERhŃl�m��^W���vǪ��rN��%�*���|(� ��e���0��3=V��Pb��Z��I�W�)�:�0h���s����1}=�:s��O<���sMT&Et��<ݱ�\�gm\+�5���c^2/e�s(BJF�Us�r+�{�5�OξXH�o?ZBB�3=P�g3�uͣyI_�xQ�y�E�L������lʯ��@��)�pAV-%7/"��ލ�1�b�:p�<s�1b���4�`ς�~39YAw���1p��v�Ր�ţ�kAa����LX �=�+jb��S>s�Z�����	�`K�e%)Y�q��_��*��!�`�U*��D�c�_��n�sq�PZ�F�NK��wtp��l떉K*����a��/]�旄F�P~}4EوňL�a~|i��fl�o�M�@O�xm����%��l�b?�����=X"�~��-�@�(~���g=)�6���ne�F.{��ͱ�ȧ�P����W[}�6]R���+��Na��2�&��<f����P�W�-q��)��*=�}��~����_�	���.�è���(ܛ؊�o	;yQ����ƛQ�%:��%�z�����QpW��
]�º�S���g�g����ί C�z�@�L%2*a&g)��W�rZia������$9
t�GFjMT���ǯ���e��Ͷ/��^��q9��棺��+�+���7h�IH5�׎�	5�h,��:%]�<��'�*e����3�+���D�>њ���>����>n�[؜�q��JL�C�}�B:$���Dp��H����u�<b��9׍vϖ�ڎ��/��d���3i�t�4r���qE�UY�+��h]���ÈM�Y<�I�,Lb�?N�u��iA�z)$�\�
6 �D="d�(��1<F��Ws��(�
�x�Û���pg����t߄��Lr���|�罊��E�M�`/^�����H��9�Ɋ���υi~#�h1i��M�����}V�d��뫶�/�[8U��(j��2('��H��"4�P�r��]Ѫ��J�:5z�0arћ���c>�ѕ��1P�Z����"^V2�����%arҭT؍�L0{�rT@�͒�^rȸ��d>c���� <�>���j�&�1r��d�ڑ�R�=����%�m�H�V��T�y����i�fڏ\���V����7��َf��7��6�'��t��"�l^�b+G1�#�(�3Ͱ �,`u�̜������RI����.UcQ�#Ԑ�p�t����J�&
��{�3���K�^g 7R\o�s��wx5���keQ���9v�p�G"�U��u���M��⌚.���r`!�ܦ�ӣ ��>toM����~�y����ͦ��>7M
�2�J�h�DbӮ ���H�_QR��o#^��85F�5ȕ:_~b9�I��
���VJKm�?Oi�5i0mF�2�Թa�u��N59!]�ҽ��^@�I�6�"��%�0Ş�;��g���0��}� �?��7�Y�/�JQ�C���e�0Z^MzyU��t���y�c��P�ѹ�xd�2F&	`�ۗ��@���]�����[a��~Z=�+�[�c�d\�f�����Q��ⓝ*��):��,Ds[Z�LY���$�����\��W1���eԢObÌ{hGk����W��ާ�~rs����J
kR\�{DP�ܜ�K(){�BRRm,���#�/�h*��7�}ɽ|&��	BE؏����`΢�&tE�S̆o�Π!!�#�氤�۳)=|x�|PY���ڢ��jd���{
��F��!��{�C���eľ�xz�x���<Ӭ�T���r�#�ǃ0!�����B� IQ�Z5k�-���N������W>�`��}.�@�6�M���ʖn��j�+T �����eޖ�����CBI#j��2��Y�A��O��C��M�~C�7q�Ct�C���~H��a��z���fO�^P8�������]+��3a��t T�O7X�|&)�hM�����?��q�Ew��v���K(|�����v����Z�K�e��w,��z�kw��SL'��r��0�p!�phH��W��e�uI���ƻ*6�`�]x�_�j� 2����p�R3��_�&��C�ކ�xG�B��P�T��u���<gs�K��tń�yتL[&1��u]f59P	����G�U�c���=`�����.)��w!��77f2�;*�s��X�1���Ŏ.�i�յB�14\I b"nb���T��e�
ԟ���c9�x�ɡbw�#у�J�|��Z_\Ѐ¥F8_�m��z��_���6���K���o�I����e��Av:��e:�%�i��,`
��_UB��?
��a]��H�x����{�#�J�Ĩ�B�l�/L#X��v��+��T��v�v.�,�q��]�.z�UF{�����b!�;���KHX�l�_�f]uMO
�b�c4Vn툥wyib�3�����m�� �>3В["��CxE3?U�� ��U(sRK:�P�A�S�RJө�AKy�C����'�89�q'3�fh�y��Ѝ�nl�I7{�OrtY�s��M�vJS�Դ%��g�Y�����h%�{����`c�!ǎT�� ��Hr��Qȩ0h����I�v���>lwQ��8��b�rV�B$#�����<�]���( ���l��}���O܉�	Yo;�v��|���|^�+\B嚍DA!nc�䷝�~�nI+f�2��������bJSB�[����gэtP��K$����Kf7�G4�i�|BF�e'�� ���
�Q���D��񐿇d�6�/�P۞@�3h_��yKB�̥
Zj��3u-���|+!�9�7^m$�נ��l��d���jkV��i����D��x,z�7�AA]��usCeO!��O%؃���0CSva��Q�`8�YB���j�Ej�)Pa��s�f�Ӟ�VM�J�Hc��'ɱ+� O�𙸸���;�;bD�RL��f�97��2{��^{�����<��x�/{��`y;l���c�	@�R�����<La>��3
�إ%�P�T��ÿ-�^����Z}ޯ~��٠r�*&�/$����Y�)�x��������XL��moD����40@����˦d©M�����c��1q��Yng,h�k��L�6�^�,�X2�l�5c��1�h��m� *�`h5[KP�z2�=]M��:}��ݘ��ep\/�󮰨V���*=U����T�vS}}�*����}7�r�Pm>l�?H�&'��[}�x�.�L�b��'��`��AvS~�*��/,�_�'��_XZ"T���W3<}yX�)�׺�����PR3ڒ�v|���jϱ'y8!�4}�c�k�E��ꮞ�&��x�$��fZ ʣ�b�MR�?�%x��g�R3�3^A1U�蛬������Zg�) 1���
�)��$�(խ����b0,���Σ`�� $�'�F0���^q�3�����s[Z��R��E��*�����9Et)Id) p���:��3ű����_��O��Pg�2�ʽ��V��׻`�cC����S[ք��eb�q�n������2�vHZ�l>�����Yf�$�0�j��~l��R��o2���)��堇Y<�]G+F`F}� �$��A�