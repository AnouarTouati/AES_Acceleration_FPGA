��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P���s�P��	�?+��+��1!�Q�u�\�yԨ�)<Q�P0��e�_��5�����-��w�t-{��+ˉ4��+o�`J�UU�s��cy�P������1�~[U��%%a�q�,�ڪ��=-�P�փ����?�O��A(O�ț���{��d���&f�ys�rZ�P?���}׳��Ĭù�c��5Q��PX���B�FW����a��/� ��q���7�*׬�������%��A�>��Q�6Q
v�Fw+�_>}^��[^:^�vDϘ����h�jN���W��.L>E���<��|�<!���%4�f�=��OZ���"��g
=fLŚ�	����`k:�)�X���'�XO/u^�ر�k؃���Z+�5�@�epфf�������@=v�x��!�4����j8sq����KݩϪϻ�\�s�q���{�R�u��"�����wֳWv��0�!sk(#R�ݚ����M�؈2�Ac��γ�71�g]�J�7�qH=���Ǯ��v1L)��֌ !{�Jݛ����0o>�)��9��Ȯ�K�,�u_������#DX��Y��V��q\��-��̊�'�&��k��� qH<^K��$gBG�vn����3	VJWKg�Uh�(�����]w<>��G�j�8�3l��%�J�Ը���Pk� n�{D� �]đS.Q�����v�8�Y9hcҹb�����']Q���x�O
 ����c��U��s��y����"�b1�s�N��g�~��E&����:���vX�U�}��J �!Rݛ��D"ԆWk���f:WWN�w>�#@\@�4�JKn6`&����3�	�Y��i�/���f���<W|T�����n��+)����>�����5��j8��,�^�NZ	�e�A�=�j�G��	먧ʯ^,��Ξ˞Ψj�.���TCk��c�,�!~&ު������H�`S��AM� �ֻ��! �x5��{�����j���C*60�5�[�^��wQ6����!��Y�%Z�}���r��R���k��_��A�v�О�C_.�t��^Vt� �$����E6��N�QQ��N�P_:�'q�J���d�	������=��p���v�&s���=�sY<�����$�yY�EA#�	��)�X�f�Ճ�,�J{��Enc��K^������+�pӻ)�R{��L�@>�sY�]e���'��y�" $�-T$BD`kx�#B�)[�Ӏ�h]���r�[�N?K\|O$X
$_�vL��s���,:$��.��)���;�W��Lib��_��fb���<uR��ML�6=�/o[�dv������2#���N�6�RPC]zk�ј������0��2a�y���ǭ]���vZ�,s�{Aۯ�����f��U�^�/� cf6��|��s��9��^&[W�:���)K��&���j<M�q�������vi`���\����3�ye���8Z^A�Ob5��IX��r]]��P�:	2�F����|�
��Ǎd���p��{���bٮ��a�=�n`H@�T��E�q�:K|��Πz��ϫn-���Kt�>A���Xn&�_t� Z�Q��
hw�p�2�;"�IQ��~�ʵ
���E�25��YS��Ҷ
���lop�D3H��:��{�oHG�W���ۻ}jw��??z�h��r�u��NG�,�t��4D�i)b-�ADR�bG8"��DM��i��Ö�3��#�^������A��L�p��sM�Ip����.��ٱ�R���og�x�s�zes��6��V�c�+�|�[a(���" �y�|�4�U�2ٽ� �a,goyfS�9y>�l�{;!v��<\�I���T~�Gl,�z9��1_�VȽ0Ws˵P�s)�A.g2���D����H�	׀l���n7��(���]>g0�f�>�!��WB�Ɵ��9LN^�垵�h	��8���S�;I�
�
�<[�Ic`���Ui�<�J�C�F�0U�.U1iI$�z���*8�cJi�{�4s��h�5k]ⴶ����f��%;m~�6/��h�婔�/j�h��az�4:/^�b����7x�q�<��������fڹ�>n��F ���#A�RE��}S�eVO ��]�vK�&jY��	��V��,���(������FH��]*�f����@�2 G�d���M��ruy����X�Q���������@.���<l�X=�H�Ԓ-X��+xT#{p#���k.V���TX^�ӗ�kDa;���;�.�w�~�1��<����KK�M�2Z�I`=Ǜu�D<�Tt�V�~��^�+�_E�)����hc�WS�s�g�������KA�3�~���x���Y4i#РK�|L�k����y��4��+n?���@�-c{
�x4�Q
"u!w.�&�,�W��3��pk��B�tI;a��6�U�Ƽ�[��//��2��Se��oB�|S5�Ŀ�y��>���u��������W/�sc
!b��dG4��&%���I�m^L�N?����[�-�jōL���i'f�Hv:m�����v�}<�?F�=�y2@�TS�������?���<�Z5��	����I�p4��u�و\�LI{�Zv�^3.p")�;����`Kx��� ���݇���M23�о���|&��Yز�B{4�롁��*�e�����ݨQ��󉔆���:�+ad*�6Ԍʊ�'Vo�{Z�������7A�|�f^�C��O�E����ΟH�Ɍ�����;\����W���l���M� `ob��R�Xf1�ԁ9��dpX3'L60R�R��a�⢙���R��+r�^��}=H�̡^w[�T^I_"���O�R��r#j�v��\����v�%l`��j? V�A(K�r��tB<$�y��u�N���ɻ>n�ze(��`w�J��3��U�V��[�{�[[�����D�B�1³���6QQ�
̸����Yy���;z��/+@��:��Ϙ,��I�]G����9�l�c�7}����^�YVs*��%7{���w&��ߺ��5P\�Qt��L�������a��s1���'�j~+��yѮe���*�r0K(
���:#H�36i����O�(�:H�K22x� �*�q6�����j�
>���5� *��rnIM�Ic�9(5��
B���D͡���A���~{V�B�1>����������y������62eC�Z͘���u����L�59~~~��,bV	+�L�d��n����]�� h��CT��h���mzBþLt����0!�sJ��?�]�^��f][��j�Ŗ!\	%l��mί	����O]Uo�4:U�
jErH�L�W����/^ 9��l�d�L.���~^J�	�����:��aQx@|<iN����?��i�P��G3���j$�W
���*�'��iNv���a���������Ec0%�~]�2@(3Z��Ǟ�_h�z8��H}��?�X[8�>~C�p��ܦb�C ���bȿ�zu?�qj�'��k6U!Za	�y��ЃbJ+&4!��`��P����->{����֣�wm����m���{>� Ѯo��e�~t�_j
����MpA�l��AJq�O'�6h���L���G<ɢ}L%����RW��e�+#�+@u7��FL�%�|b	��X%�5�t+���-�ĢY߿�O���K�:�η�?��|�6����c�-!���Iχ�L�Y�� �7�Rw������q$���NcUȁѸ�"��;l3�:3�5���V����/OA׷�����-�mВK��.GRE����AN ?z�I�Xk�CF���nB��[I$�e���s�3�>Q�@�\2g�&�{�%�`i��S1�<q�>��U��!�Fp5E��^��K\����>��;�v��ci)�Lޕa32�,�-�T�H�.��^z�V���=C>@�ʶ$ZM$٣��M�����H�D�7�5���@�_m�z��7R-�Z.�������Dg�Γ�L�`P�����ց39 "r�lM�������>F]�t��;�������G��:T�"y}k͑�fx)"�h�����J��-5N󟢡���&|�"��Ĵ�ռ�D'�"����@�qSaI���B���l����~w�Ձ�)]�r���|dˇ,���'�}2̇Ѩ
J�p���oiK曐��(��m)��dĜ�o�h��!�s��E��X#ﾲ�B_]���[�V�.�C{�om!�{��E��y��E�@v}��~AP��mT��lWL�E�{�@��<&��7���XO���� ���ry�H��+���S��Q����!�~i��]����
$g�l_���?-��RŔ��U�xʸ⪑�E���։U�=�/�En3ow���f!x��骟��c((8=Ť��)�;�8ޕ�"������0�*���b�g�G��Q<��d5�c~���b����F:`V�*W��w{����X�E*�>��R(3N ߧ�d��d�<D7�;yP�/���CS�k���vy��8�Q؄�*��R���y�R���mAԲwlvań��/)�K9ː���et��P�fM��.m;0_QQ̬z����A�cZ
_�k뱫		
}h�g��a uJ�DB~D���T�&�K��p(0h�>���y������@��������Lz|�,Ps�m�4����}c�S�̚��J��� �����!��n^��7���/f�yD+��� I������(�T��&׍
$��X��Ey�RE)��+ϨpѨ����/	�fUd��伩�u�P���Y\��1K|"7�d������L���Lѥ��go9��/Z{�T��C��d~F���8���b0}v��Н"��b�^���Ȟ����m�>��e����3�V���$0IVۨ&|��>�J7f"��#��C;v�������c?I�E�k~�����i� .��WԬ�}� J���ngD���Z��'��C-��|MIw�D��F�Ů��~Koh�vo���rq-������.�įmS�Ex�q�N�O��fa���[y��]Ɨd��0t�����ҍ�Wt4-_�[t��u����`�.���}��Ew�e�t�Lz�,\x����8d� $��`�y��>a��[ �]�yE����+��v�e���c����uZ��w���À���><o�q.�B��W�B��*H|��Y������lXṋD�ĝl�{Tp6��kV���h�%i� �x|2U��Vwt��I�����x�3�`�	������>��ԧT�#*Z���c�i`���Ճ*ǹ��4��:�A>�?�k�-/��w�����`�1"�L�&�!�R��$lˠնs	��n�� W��QQ8�wBd��_@� �Pz��;��n�M<_���4p�X����A��}8��y��[�� ����h1�MX3�U#�d��(�6����Љ&� זbx�iP���Ω\�f <tE�HN�k���!�q5�}=4��U���j2��j���h�lN�d�ġ�(��[�9�BNN�R�`�&�#��lL,A��D�S# cB6hG0.ʻ�=I}� �ls�,<4B�ΐ_u\�;7�?������X]L��Lv "3�z �3������\�F�¢�����륲�]�m%��6��sz��#>n�]�@~��8����s�~�I��a�8��:�0fg���+���ߔ7j�EBZ�L�h�^��}\�nd�"�qΚ�`��L�����@B�j;7y�}��غp�0]�6�# r �?�l-�z`�AUz��	����@�?y)V?J奻��R�E)�� C0��H�$k��\Ӿ��{�$u{�a����![���c����g�2�]�͌�8�!�z({jHl%|��7q�z@ᱹ�fx�� ��8�J�*�>?�	%��0���^jDs(�,!
9��S���kÓ~�=�j�"�s)���8�<{��:�\��~H�p���.�Upv0a�(FE-��ݧ�Km���A��TQ��cY�q-����>#�L����T�`�\c�&Sh��E�������wk}�U�	kk�������;��@��?�?٦m�\V�l�4��V�jغ�*����W|ӄ�	�ڽ�U�8X�ŕ&|\�|lD_�:�%���r�cM�9�_��L��Ӷ��Ӛ��﷊w�Yu�4�o9�$J����q@���@fs}���p�p�X�A���#�w��/��W��NMl��@JU,�=�x�W�#y8>��+���G}R杝;n�������r�)Al=����T-�;��739�U�P6O݋���_�u�<ړ躣��hS��H��ćߑf����G!�Z���'rK7��_��Y%ߤ�X6X�k�&ζ���j.-"Z�!۞�5�WC��H�b�L3�
�)�!2��9x��3�^���۸���N�����q	!��R�������SA�/O3ԙ,����V���Ҙ�:!t���� ��3x[���%��~���;_��*�o�L��u�DmL�9:Ok$udp�Sݍ��n�KE�h�7�>��-����H��Û���y��}8�/CGvcvOJ0����P��ݔ��0Ͱ->GO��I�\l��P���:PNR�{��@�0��B�X�wg����x�H
p��Q$�܅)�(�/l�稩��`wG"�>�~��~{��yc·M�"�n���F9�����#��0��ß��/*f㳪Xr��b�n �j�R�{��f� 6T���|��Ί�P�|R���������-�E�`\EX���uC�<><��~D��p�u���L�~X�����~j=��?\����Ǌ@IT�*�@��u>��%��&-%��Y�O����}�L"� h��LNj���^�7�1;�A�&V�	M���5߶ �Ѐm���2��`����A٫���ʈ,dټj�Oc�ܟ�+��Bia���Wq��ä���,���7�C6�{ʃ��!����:yF\�]4D���qݔϐ뗳n�B#c� ��5���8\�f)lV�1�X.���칷9͟����P���E�Ϋz$p"���:�W��d��
�SqG?Te���l���\�~�Aw.���l��������g�.l�Y��I|>��k5Ѱ��|aχw�5-���Dn���!�W��P��^���!үq���'���/@���:6��4�𬔞�BH'���&gj��;�.�5�6���#r�)苸jI4G��d�ց\�5�H"�T�i��ۀW�u�ǡ4q���oCL8���6?������i�+��Y/'��Ѕ�m?e��|5��'�j���t�������"R�5<4�l���{Hu�Is�Z6��W5�Q�t������5A��7���d&9����H$��c]��|�{�������t��&�<Ŀ�l`_R
,���E
�����X�1Љ�Fm)'����4G,iA������$ʇ���w{��xs�3Z�����Du�	��o�7��q:1RxG��GҶBu�q\Or��/�&9Z��jm^BW���}Bk��5�ER� ��¨e�x�˩�����d/:�C���M)K�T�M'�~i�.�߻�JA����.Z%o���Kט�)�-��2�ޢe�H웽$���#�ȓM��ZLc�㸞p�#f���w��| ���Մ�*9h�dV�S�6�Q�n�Qu��k�_71���TT�Ò�|�n��K�G
��Jnؤ&�`��CK:������c�u(�g�������]��}#�������3>�Qc�Iꋠ�*�"�(�U�WA�����y)��E���x�y����I1�M=c-j�42��v�܄�s���������}�VB��6��Ł�M���vT�=k�� ���_y����u�]�6X��������V��Kke� �4���{�R���h�@V�	w���J�P-�Oǔ�|
��X���3,}Ims������UT��Ϥ�M��8�t,��]��+4��EԱU��=��Bp��d@��r��ՙ8 �ۍ�rK�h�2R�H9���,��FXL}	�#TN���6_v��k�n��z�`l�>�ѧh$��^����Jo� ��	G�8J����.��F�с�θ�Dbr����/�w�lw����w^��HM�؆�&��r7w��I�޷P��G�y���zj��־N��Y�n"�sy-,Ͻ����	�χ9 �*���]o	l���+GqI&̄�ʙ�@ѫ�DL����}�^��۩�5%-�V!U&�u/�|�c��_��GQ�̐�,#J���õ�LU�^�9d�.�ea&��:��rM�$�;�%��"2�F���S��"���(�����Zh�_啰Y#�;E\�B�l�N��Ȍ�Go����u�T�[q�.����M�OMa��Iߧ��{d�c��ө�)p]DÙz�+o�v�sH=�Q`���HE�\���FB�9��K�<_�#ms'�Ç�km�K���L�*���1~�]��cX�Ep��W:p���'A����c2;�x�E�
����E�]2E`�:g�0���/_�N���!�k�!;�2���ĈN%U�E�67E��fMIp��bD5	2Ơ��
���K4g��7|(e�-]l6�CoS���]H�"!��X׀�/ܬN�u}���L+���ݬ��8��CuYud֊���E1aF�+��Ƹ|}��j��Z�ץ�ax��W�	1?���!Z�.�~�����|D�ɨ���;�h�D4�?����p�k�U&�V�����N=����Z�:��'�L}�	u�������|4X��~o�v���n���C�{�j`j`'�_����#BlڍԦRW7v��9��~�� �t��@�ʐIK=z� ���=2�����fuƀD�:��/�G2W 2h�VֿB�=+�`�����<�|��(���t8�c�X�z��&�ͽ��I�F�9����+P�!ɉ&���iwjGĮ18Ren�nֿ���B�Ձ���y�vJ���1��j�rޮRS[wTo]x�HM��qV��*Ջ�Dw�zd�t�:�B9	�~l�lּre�� e+F��~�//��+���cH Vس�Fmã���hg΁�g����]_�9\���*�@�-:��A.�J�U��n:�if�]�؍�7�s64DNQ�y�S8d�j'�א�]�P��m���U>�9-x��zi�ʃLۉR�ь�λ7ofmp5y��+��B�7k4=r��{T�yn�Μ�3)�T�O1��Δ8N����87qM���K*���AM��q��>�	�iP�÷T-� r�΄������{��)�R��H�о�e�~v��izz�ȷ�J�~=�>2[(�y4��k�-��*��t�d?���@�an��bq��I��G�PT�����I|fy��H[yGb �(�:�jJv��z)�� Y ��I� �
�����<?�-tػ`�%]�>66u�SoAF@B�G�1G��&�h�'{r#��J����"���^���>�ȑGu�<���y��ʶ�BxO�y�as]7�T�<Ș�^��ܾ�G5�-��f�֌tA��&�'�����-���A������`
^��k�ܠ���������[�Q���ͮ���_�9��jʖΦ9� ������ y��h���a�Zͬ���N���y�W�T�/ �,a�/êIk�\@	P_�qw��	��Q���U+;m�T�����Χ��f	$YBצ�� �j�B��`�)#Zq����
%�n�,U��W|o�N�T�=+Q銩����v�{���=]�wd��.�xب���l�T="�?�ED�o�;7;�n����U\���P���7A�>�z�v0�������Kh�YN�;� ��7O{H,����0R^N�)�:�l�m0�Pp+?��)����	)c��v��m�M~��"J��ls���!�l�A�Ĉ�4ח1D"N�`����0a��pUλ�?�{��
v�����D�S�0�Gj��ڂi�(��I���2"ȥ�,��b��w���n����Ö��'@�h*;c��6-��+�Z�\\���2�b��QSo�7�{��������{/ց9q	C*H�dw�r�ru�N�Ov	�I-���;�/|ńd���e|����$+8�ERrD&�'�*
�����'�� i߃*cu�M��>��HqڼZ����{���m���[���6UW�g��X�
;�ǃ�?�#g�(,��D?h�٣!E���W'a�XS<�=c.r��ԞW�T�P�M,J]�	w3���`� g��T�7΂�#�h�O_�qJ.�D4�bM��s��UF��_A�~E���|i�o��Oe�g���R$����.d�z��U��}�M�0��|�_�q��������9%���	hg�mye���WD�<�)�im`$E8�j,�G6�+w����R�K44�,EWH�F���l}�4v;:�"M��O��
��Hم�tb�#zN��Ayd|��1/V��W�0�U����3Pp�;����o��ʓ�����At�
Ջ!g��G�&�,�/�䙅�;+)o��u�Z�&1���R�1w��M`���mkp
���U�?4��q��
���w LNA֊p�7�"HS�G#N���wg�'t{sry�0ж�]I��`�]h��e�i�`���%��Z�l�.�c��s`bǆ��Q�u��
	��m�2�2Q<��������%L�g��4��3��ˊ�\E�A[r��j�p�Jםԓ��7�B��##n٪�v.0qY�o�D} ����bm����������Ksͳ8�u��s�k?�S|�����1��3
*.������E�����@$]{����t�Z�;+��6�K�8 �C<���	'��_�B[��������\2��Z��(�	?�u��͹�&�8:�Ω�e�4�1�m�m�֗�+n��T���� �q�_�O�gپ&��8���I�HJ�ZZz���6f����q>�)��~g�!�����V�֤�J� ����}��lB'�s$��~��	��i~��pS`�c�^�BgBs�|^<�}�Ɍ���5>�5�:��zj��pd5�+���jG���Si�E�<k��Y&�WO�_�2�pc�b=��n[�P<P�	sA��OW5�p<W;ª�A�-o\}w]�+�.�%;��S�*�jg�ȽYW�SHR�vN�2cP�]��~u��q�0R[8D�r���.B����[�œ�!Vm:�&��o�YDc�D�Z�r��1����kjd(��o֡c�/��i^ibT͌�����qLx������UzL�N�n� {�!ĴUԍg+����_
��7�*�'��=�w�m�����%3R`���+e�g8t>�˄�D���~��m4L	jf��
k���rW{�"�Pd�H�)�op�O=�TӃk��a��SH���,�=�`(�d�62������ࢻ��"P"Zfˏ�����W�Qؾ�,A-�=`��8������m�~Pbȓ���i�� p���~p� T"�Kg;`�ڼ�Ρ���f�ڧX�<_>��V�@#��'�k���Pn�K�p?9��w3O&G��^$�(짃E-�^�d����P�Rf�p�uT�	 �?�C�t(�C�!�<m�0b��6s�(|=_&���O��}���D���ٗ*����6������v����|x�dyƁ���u��/�B2$�6%��V$��S$��t����uV�7�c�f�0��t�U*	��vg�������\�&�|ճ�>͒�E�+8�]���W���]�U0�c_��Z����h�1]J��g����2���3 �b��"�c�~��F�u�sk�R�O^]Z7�VND������I|\�s�#^2vOI	Ir��\+��A�!sѠ�ܖ/�3VN���N~�MS��9��i!�D�iٴ��n�q�=+�7:ح�U�Ѐ,NǙ�5�e3�8i6�7)J�颱Hr���[��b�p��2�pO�
���.¨3��ᓆ\7�MY�����?��J���~r�Y��.�>�LH���Bo�ɶ�hE�����c�ɐ�u#�8���1ZR���܍Y����TcCI8
�*�x�gK���=!�eڞ��ޛ�//�fL?�����X�#�I���q��[�
��T��3��W�X�h���&�����i����d��b�68�N�E�εL���'XV��~)�[W(�g���,��>�s.�S�dO�U���ђA�B���i��LU�vy�!Q�����Dj�3�1��5�-��RסS��lQ�����ޙ�c��l.&��e�k���E����YU��my� �F�(�0H��k��ǙX�5"xG>�ϋ��y~�Q�\���N���p&@b���Q4r����4-��QDK��$��q�R'��.�� ��/�
���x��z � TӠN����D��&���{�\9�����q�M����ͷ�Л*4t���'�o8��Ö��f`i��3�r^��/ĕr��B���������&��]+@�Ԛ�����%-f����y ]G�S�fw����-�J����&���oũg��M�	������<��t�s�e�^�@5w(��Z̰$����M�R�H�
��,7��6=#RG�\��3v�X����p��G)��*���&O�!�����l6�\��G{qHW�6��9�H���z�IK���׈3G�����,����;U�^���ˠCTE�x-Lvs�Ӡ�����D[t�����NA���/�`�w��5�6��/�V�8Qz��\\��	Ik�*�=��k=�"���4�����y7�+�z$A	²�l�}X�r;ɋ-_��	7]bEZ,�u$��~Hy�w�\Ji1+0�^�����A'�
��c���}Tjr}B\�~A��̂��m�K�W�5��p��Ѣ�K�=�����&��t���Tr�Tl���a���݁t�G[�.O4�]F\�E�En��f�jO���Kr<��$���.0Q�~x �3�NԔ���K���"��/���A�+�s,"���Mo�j��z衧H���J��B8�eD/v��4�� �gap�87�/UV.����Iy��T�|�J��i�a�z�:J�n�<��VD����
�h�.�Eh���?��r�p_x<��o���Z2B�5#iu��M8�=��ڬ�����6K���'P#*�B&�5���OB.vqA�kT�NF�u�"���pWA��cUފ�l�ˠs��T�g�,?�B�|�Ȃ@��!:E��R7�z)�����?V�D����[��1XLd:�S��:�0G������V��q9��P��b��<������:�(
�KPe��z�(w��ݸ���p�z�E=�y;e2{�R�%�퇡�\<yu
��V�p�wR��,Y��z�9��DGKJ�R��v߹lħd]k�o��	��X�i��Y���0�r
���|��rE��y-�y�d�h�˵��b�y	��r)���E�͸=q����}�~yL�2v�:klv>���F�O�b�(�G���<��`�o�^��Ŕ" �v�GD���L��$:��v��Rn�k&�*\�e��W��@%�����nB��[׎��b,?�\�&m��8������|+��D��=����2�k�{+a���p�j)�s�:��"e<��0�E�~�~�@��:E}�H����HT��.��fa�׃����ZY��64:��A��8fC��!ب�xoc1v�h&?G��?����{��4���%�3s}�J0<��z�'���m���t�e��r�zBlbf�g���铲�^���u�i���<�۱Oփ�X�\s:�Nbi*��d����ul^4��jDa�
p��2�0��=�S&v0�������!�
�Zq�>�L��(�?�.���Y�(k\�r�>��|5���w��eԍ�q��%q�x���P��L�l�KVٟ����s!Nl����w�t\b�2�A7�޶�;�U�|��w�R�6 �,O\�r¹F��cWY?Yo,�w�_nk��l�R1��%8^���r�M@���)��*=yc�+�:�"Ѿ�4�6���/1�yO
l�<[&1;�
@�6ݥXE���ꜙN�U���u0�d9�X��;Eh��h��]V�:ؔ}B"K'/AN�AL@����xS&�����nE?�l*6f3��*��ŀ~��L8��3�+��[�>@=��3��%�d0�\��W��lW9p���,/+�@UIXM;�Z�%;���)�L'�ľ	��̞�-��X���G'���绝�Ģ����d�U��J/�t��Xl4vl3��5��v����~%��'���8W{(y����0�81�k���θ�Bt3G��=kT��u��g�F�$#\�6�����tB&e���u�*���e����o�X�!��MZ�'���{
�k��A�h���"��?3�/�4��qk�}��"��(��
��N��Ւ�7J<T�b�^�%~4��4II=�|��ҊPl���W���Du&������{��pO��G|1LE@��&�:��q-��&���9�ٚe�{/h�S/К����{�:��O��j��k��@$"�iOR����Ω����2��˻��K��hM�==���A&�K~?N�c���--�y��j0V���Ufb����@ �A���n7�����@�GV�ێ;��5�<��r��P�ub@���&|H�J������u�b^�s:L���o�2���|���6�"��r
M�O�)���ưA���GJ~���� )�M�wE;C��-����O8F1B�RI�C>����av(��/�]64X�����.���e)|�B�_e����&Tl���R&`*#H�ަ���^���=�9�14�j�O�ކ��V+e@�r	>�ꉎ��u�P�'$�
>��线-Z�-'?#q�Y�ߤ+�U��y�$>/��B��X�a�+i�l��e��g�Տ���,�AG���q|܉%帬d��9-�P�PT��t}�D4��4�6�!$d��.�ⴁ7)RzEv-a4��������QwS�Z��ap0i��\�%o��{]~�D��J1�9��p���t��OJ���
J7٘�8`|�D:_��_��8�9�wfL�p��J�wY莼��ߑ�x��i���7�"���d}��9��?ܨ60�pN�������%5x��]�<8��QĪ6�?�8v,ί���Ѫ�ʣ1��<�����'f�~�zF��(���c������Q���Z7��_�����6нχ�85�ںB/c@8>�P1��q��&0��U�M�ʱ0P�o��͸Z����~� 3�ۢ�a(85è� Jt"���O�����l��N>���>�!�'׾D)�5(@17{������5�
�wر�l�IC%���9�&{2B��z/klǮ
�����F;�3_��t���Z���Hv���5��,���9b�qD�u�kА�-@㌽E|�	����fOD +�91;x�o����սo����KsI)������������|+*�8�����X6�u̟���Es�7=�r�����m�~���|'�|LE(|Q���f�#g'�R˃q}�+�/�0$_SD����ca=>k�M����}Ξ��R��9I�"o��mY�Z��v�[8��6*�c�gS�gl{<��8�u�G�t@�EQ���^�OY������y��*�U�`:j�p�N�y�u�P���Ԩ�9��7��@X���J%TՉ1m�7���?�6����P+� Q&�ժj������,�؍����E�f"0�%_-��󵚌栎�\,`m(}�3<$�pz!��|
��}�����N����2������0�
�E��s�����J���C[	`�y)���J��K0���R$�unl��[��|N��d�� YO�fɳ�L2Ѩ7��w��D#�Ò*p�m,㝽�`�(���D�?��8��ky�e�Yhj4	a	�/qUeH��Oc�(j&$�؊p�ω�
Q�3��
�Jb��[vC�Ϟ�[�w�e�3k6pwl���VcZ���Q�����x��f&�d����i���՜�d4 �y�l_? "�01�lU���V����ی.��g��GWAN��g�3�s.z��> ���/���s_M~�ă��
A�",�IO��נS�JS�� ����f3{f�ɋw�<dU1����:���^d-���ʇx緱��������Aa���Xq�������	��d�!��ċ sK]����#��F��+�f�UE�h�~��sY4,�T���(��2	C����W�=u8�ߌϊ�Ҷ��s�U�2�3�ٚ�*�:�?��OG%�a�]~��{D�/o���N�_T߈���FW��Hr��n�}���t����s�H��onHC�����u��Ӡ$;r!���[ � �h3һe(*
��Kiǝ��m^�p=�|kg�~��c,�b�md79���19}��_����/�@�	g�OϚ:��9Ѿy���Eq��`�	���k����?�P�<���k����K�G,�m �ũ���r�疌���E�u��_�W���bg�;���逧����`���W�A���is?֒i��T�Xg>n����������ZIr���٣�4Gqn���r�����U�U̯�cxw+�k��!hK�����p���0�#�f�Sd����j
IQ��`��9z��9���yf���A�
xDC���)GJ���T���0.Ð;ʗ,�*A`�f��"d�����Z=gcj952�4���<Fw�����s����hbRs8����)��j����s�i�	C+��V�SU�5
L+|GB_�Fs�1��I���8C���y9}p-�RE��u����(��փ�/=�1*aN�^g/��f��j�[w���Vr�6HHq�w ��&�Ҥa�HU�8cXa���a$rpW#��&SjHK�;)Y��!'3�B���٤��$��>������P���c��IKzX@�v���ʨ����XkԘ��dǢ��2�v���z{��Q �A�X4����A[L��b��B���ߋEJ6Ns�ID�cX[��d��E��eN�#�"�|�d��	@��&����elOs]��&�Y%�e�j��E��Sj���o��~s���/p�6��Iǫ��z	]M��4A�;�~�6�6o�-̳L���ڇ��n&D���R�<>��-X|��Z�7�[=�����>�oOy �n�+��v&���
��N����Y#�`�ߚN������^�Z��z"L'�������#�Ox�ED�a	�\�[���X{���h_�K �~� �TZ���X+x���;�?���R6_;�<� ���	[���J��q8")�G^7�|���剦�++�����Ư{��u
���&���R����K�~[�i�'
)@HF�/��o���@!Q���l�T���P(%v8�i�}��e�ú�H�O�/'�Y���wr�4�uS}"d������	��g�F�Z�X�P�_!�W�AmC�z�m���ٗ��!�-������6�s ��@aZK3H�1N�=H�c.ԩ�̉�E.ȵ��\���;��TC�)�*6(��xA��M'������!��T}J��jl���K�+Hxr�/���IZ�ź�y@Z�����>zCE�L!��uEcf~LTE��I���=F:RVO��Nu�V:HS�!xC�/�?�gS�\Ua�P��"	�z�u�h��}-D4'@V1���E������$萧m�*��[��<d*�U�poʂ^�D������=S+�f�_�1�v�j���j�(��V����t7�ڢ )P�X�fm��4Pox��	����&�V�'O�R[��㻄�mϚ"im'�����H�,�G�EmG�t
N���\sGc��>�3�������ׅ��"2�m�{�����V|��n���%۳�WN���
@��v��U��&-�&�o�?}�F&lYy�+%��E$�}���Vu�'��(/ǡ���%��
�d�J)����W� ��^1gO���֦1�.7�vv/�q4sa4p�Y�,�����t�S�[s�����d �7�x"MyW�������-!��\�~�����Qs����&+��g��8MJIY2q_�ړ^�DOdOz�Z�jn}c|+ &���^��s~<�������y�w�u/	�C ;�^G(0�Y�Nf˥��:�f�W����O�8��j١���z �_谤�����)�:VE�
=b�Kf��yoT��1{>���$dsQ:r�����ˀs|��Y���S�����M���#���m��-��(]F6����4B��:\�]h}��H�'H�����7��q2	gf�4����q;�ݲvC�\%Yu0u%��+G`���~�^������J���F�� ��3�՞EԀus��w���k%m�o�IA�8�M�����eD����I_� ����w�(�x�eU�,���Z;aW�yd�#���K�aѳ�lU��(���KS�u����8'U.&�S�WTsk�Js��݄^�j���>�`��zc��4��X@F| ��
-���y�GoD�x=xp�p��K.m�?�gP�L	F��k� ��YFUb@��W�=b���X �0�`��.,��8���؁IQ�-�����-����!�r���=$��O�vJq���D���W\"z�4R���|X���LV��}e���nl�*ElEba
�w8h,0�%-�%o���������߲?��EA�K � Y��i�I�s�n�'��n���,�vS�bT���dD���e��p^��Y{9��U�e��A�ٕDe�f:����l�%��QI��[Os�$��:�ٳLe����4��m�۬^b6�=�UE �U*��jE��{���#����y��@�r�u�eռ��,��ߡ9�gd�B:�V�&V��r�As�Z�/(Y���~%D
��tR6�Lמ�c��O�N�7����y�@.�+��*���r�
���a�3��"��`�̀���4 ۥ���`)�k��1fo�mQY6��^�x��ч�}�L�������[�r`1M�a��ݼ����'P��L��"ˁl��t��-I����B;"����~G[�3��)�{N�"P�umM]�1?qd��$� �5�u����&���e��5sh��=g!CIt��pWюk7�%����M3k�[��Ĥ`AI#�[��+�����+�"�e'�s�� �޴(�h�����.O���V=���{l ���yؿ���Nh�P��W��	�h/1�z�.�����sh��?S�����I� si-���M�/ӷ�=�"G˗�C��T�N�b|�"YI���d�Y��I&4#��ھ�}DX�}������ۗZ(S�-�LK�@{�/@�����Y�����zM�x>�"w�!�#*�M�n*VI��> a�������0�p�zQ�7���.,�TDͬh�>i����Z��a�� ����Ɠ�Z��k�3@(d:�>��x	|h�м�5B�����	�����nָ/>D�6��m�E$�%�BD [����Z����NrXV�z����xFA�n%i�2��]f��Jl�a?5�5�O�T/��%�%z��z��ձ��	�������l�4�YN����,����Ʉ737&����&�z�]=m�#�W�w2�w� ��ٽ�0U��ҙ�n2�<%\\5��|�F���Wrv$��#�O}�SFm�UDy�ǩ�4RSi���{	��M�ڭ6�wV�pJK��=jz��ڟ7�\����V�G"��AuBR5���F��ro�I��ǙXV+m��2������X�����1X����6xX+L�e��{�ly���m���~��V��������b܌:e���
$�~�L��Zk�2�'�A�jj�៛�b�d�r�O�ZLºj@�0�%{�a���VY���kãg�@�[�V4(}>9��PL�G.���rl�����؉	�LuH����L���������[�B���Y��5��C.9.@��l"��ܸڭ�}��� ��Ej��:vgs2g7V��=��]��	6��%�5�% ��<��KA?Q�&�2�%(��Ok�ش"�$�%��9� \�jC�m�ԡ��锇��M��h�c��
> �<#�N�ż)Z�Y��B��(�5"I �n��b����9~[L.�sgHy����v�a���ȫ���U�R ���]�ؗ��}�r�0e��m��;�g�|��՘ڼ>W�8O��r��#��r�#�ܩ�mZ�h��69������\�U�J$�x�o�{�7��h>M�	J�>84E�X��JI��\,�P�	@�{�T`R�W��Q��� d
�RA�-f�k\@1=���g����k�� �MK�5�a����N;F��mQą�.�!_-���f����n�òk���^FX��Br�J�ĸ8s~�Y��d�-'���JC�p��`B`3����'Ⱦ�F���$�(Y�L��0~�D�� �d�1��P`�g$?u�%�$[��Z�Z�p!��8�+�wt�b΀�C�L_�Gj��Ɨ�c$G�2X��Bp�u��4#H�L�hd���E��sm��5罒�����0���"�6�N$
�5�~�6��0��T��p�AS��^���G�L`*�a ��9.�~"�$owo=G������d�ڭa���}I�C7�����׬j�B�\p�$8jտ��5��K( Ef�|���A��ß��`du�3��Q^�pRba��4rD�s�vJ�=��������0A��Y��JA���IAm�<v~� 8L�*J0���7u��pW��b�q<�ፆ�~6ß���3Rh�0��>�`�g����g�:.C�M��*R@;�4��@z�Gt�!�־2u0�� j�[��z�C+:=�=��v<��#��$ >�-.ɸDQ��y�dA�
#�8�O�#,����b
z���
�:D,�5 �m��Z]�=�Ķ��f���5����F/�l1�/���u���� �W�Nը�(�|�i��n��邻�O�k��T������q%}A�[gH�����`?K�.����Nt�9�]��3�F������!�+�ԁ��:o Z�S��,�/�����P�
����QM6Ѵ}���|5�H�a�RX��?�������E���`dE��L�"T��س^5f^�m�H"x�����D�6q�5�ok�ц6�&��'��~ò^�f�|I����J�=c��9V�:p��B�w�)5�A���A9~4E՞Ȉ>tH2�`�� ƣ���Sq�v�'����7\SS
�J�@���E�-��Z�e��
V[�
Dli��1s�Á��^�\�r���N��(3�S'Ldsx��Q+�^����.�B�
q�����:���Z"
��jh���7���3P�@Eky�窨: Hg^ER9���*����Tt�RY��q%�<��=�jw[�����2�Wk�5���C�[tlhD�4 ��2q�!i�Ȇ�/]R?F�!mcF������E1|�y���r��|:o%Ɵ��q��
 �@��ܤ��m8=��J��?�"$8�$�0�X�8W��<u�gk��=X���l]PxPq���4}�?]��n���cko�R�<:�B�~w�JޔE�>�̎�F�2*�TWM��ġ�-.�I��tx6�A#�������фwj�J�;��:Ry��M��Z#�����2N#2�$�
{��vͳ��/�%����.;��*�?��%/�t�ҡc8��'9b�9جX]�� �#�`�llD7K�`��,O�tI�[�T���X
�����s�J0�uߌ�ʄd>,�BX`�e�! ���yuX�ui9l4��z�O��K�+BlcPfJK����@�x��X��N^W���/yi��@r�!{�=����܃
!��LIӞX�=2����G�U�g��TJg���m����B�GJx� �)M��qŘ�\Z� ����(�_��b���bǠ2;�k�G�XX=�����r����c��g�Gq1W���u}�	�Iߨ�k���h��-�����f�,���i�s����z.�8����I&��S	����qK�A��6�Nn����)��7�ɬ�Y���p�uy\���Q�ƓF�≟�ʑx`�����(�*2�/�;d�_����u��
Ri�sG���R�8l��=)�QS��4��Č�P�n����� 7c��(��L������j�/��qX�����<w�<;HUw�s�q��d|]vR^�o��k�s�Enf��m%la���r<;�V��;a,_[���o������=ʚ�5�`CV���C*�6�J�G~�x��!(�+����<�(�cM �;�jLI@|ogD�=W��m>f\�KQ���/�>*&��Φ֤r��Y+-�'1S�:��X��&%�ʀ�=;J�B�w`�Ə�eA̭,.3���P4,�6�"�y�oI�ZS��|�hw�=U�Q��(�n�4lb�rϸ?Տ��x�Nk���1����&�OBA�g8�%,�����'KL��S��y���=��q�
�vnK+;:<���l~'��ـM@��Y�S��"���QO���G6>�� �ѝ��`�"ʅ��XA���Nu!��Lr0D��N��伣��/�S�EZ2M����g��� J�D(4]�c4�)[��;9Xeе��&oXjؚ(x#�n��vD�~��ӻ�����%����r���dbjb�e�)��l����B��l�Z��$��uJ��n��~������{�Cco�����*��":�S�tb��V+&��,*F�DS�(��ab�ӝ�f��7�2 m�:��%�<� o3��)��z�^"�[��c��L�C�> WA�� �P������h%��l�Z��m��C���a��&}�rCNd?�A����x+Ka߭���ޢ�ũ�w�݂L��htc`��ա�I�HY��Re`�΄�6�B���ː3n�b��>��I�� ��ڐÆ��쪆*�E	�W���ױK�sS~DƧ�b�7���Vp#:�Ϫ��j�k�h8�W�� ��V�>�f��t���<��K}�,�4���N�F��b����H��t����~��[��B�n��ܬȲ��ц�9��YT��v ��'i�}�7���N�����l�6��@��`����⹔��oq	��(�xY�tu�Nug>�-��N!��ɒE�JX����5�d-S��U��j��7fh�J2�_S�"������q��T�4��T��2��4L�^zm�z��F�^D���G6a�g��49\ݹCx�ّ�V_V�8Vi�ܵ���IS�E�5�;�\��W6O׸t�Y56yI�E.ߧ��J��R�{-�D��C���'=�|����Y�Mk��	���p�ܱ�^D�:��r8y��\@o[�i�����	��� l��¥�!(�&M��沏n��P\3���i�������&�@f[Wh\⻭�)l�$�T��.r��y�`#B��h�T��QU��)�2���J�k����ӌk"�5O��/+~]��2�����Պ�:3��^o�}R]z���|=�,p���_X?#�!K�ު��!x6Fe����5����)�����wY�~8eD�pR�z;��hE:�ʲw�4����& �d�g{e܄�����d�b��¬��&W�I��=1�7�q�Y���i=t l����Բ�`����q��3����~]|�f�T��r"��Cr�B��)�NJ9)cPB�"�D��������|0���Je�˩��V��)��6�x���Y��&I���<��=W#P�bZ�j�`����ޒ�8�˂� �ڡ�|zO��[[[�?����r �O�K�v�t�V|�9�2֨e�[�I]$3Y[	�j̒��l�݃jv�@��g?��r��8|M�G�\�C������D���`�WG�!ua��<�7�5��rIj��'u=��R�ʎ���b��Z�r$�7cз�4�`)ㅜ�~*Eji�{���v�9�Q�5,�[��TV�e~We��Z���ɀ|�����5�*�jq��L�c+p�!}���pN [�����cJQ�-5~]Z����5��}ȑ�7+��Qj���\sА�(���V~��*r��Ñ;PZ\SܠeN�nn�N�잛Gd:���Ɠ�R�3C3ƻ�y��%aJE~;^$����ev�
C�m�IؕLi�����,�/N�̧"����w�"Imf5�+T
�g{� Ϧ���s�r��~�Ot�!��w$�l�|��r�m_|Y�D`�5k�U#��G^/�,��32I	��ZtE U���,�4���\W�G

��98.j1�EЄ�,��3O��;�rH@h��[=%���d�B�1��=�V:�iy��������,�m#Ź||*���#U �pn^�3TL�W���%D�s�z}�w�I����+�گ���X ����!��A�mrJ*�����+c�}!TO�5��6V.]b.3s_�`O��A�S�~\��L!B������~E&�;��qB�6��R�意�Ù�q������K��h~�)���v��wC��E�zֆ����+(�F3O9B>AF@�?W��E� T~����yY�,�Q�?�y�}U�/w��Ҭ��%�{!A�*��Ơ���{j�ʷB��-@%�I��P�#���
�p�=����������~u�e!XO�)��nJ����qRi�6'^�����G�d�R�]�ԍ�y��l����#j�aĔQ�|��a.��C/�)�R4�JJ^�Txf�N먝��NǷ'��h������  ���}��\M%>l���p��]M[׺��D���N�����,P��i�%9���˕<:@�:�c��&��/ ����=��#hYL�/L3���A�-�j�t:����q�I:��`:YsQ�s��G��}q��"���������)�m�~(��O�>탗���u��p�o��=��|�[�{��쥒 �����|��x�̱�_K��
�!Z��oya��Q��>�*J,r���
��x�`�O������&!��X����5�O��U�G�_S���Mctud��%�$y��?��S�;��&�$�����1�P�	�v��[ʶ�֤Ȳ�=*����@�N*5���E�5�[i�6"[rI�BI��>���ǐ^�z&����n������N�t����}l�&_)����;��^�� y��.�;�i�Cx��MX�Iy4\�k/"	,��|qq�~�E����uZ������J��a�������n�Cãh�0t�)�pQ�aA��/�y���PY���\�M�ҽܓ���J�s�Y���Ԍ�B&2i�'�ŝ��T3G��^NFC�pt�3P����X~�>����'����9��0��6����z�����X�ӈ)�9��p_����x�ɽ[ڻR�al0�t҃Z�����uq�_��]�~~�#��!tly
%V�-1��fM^�	^}TyrY ��>� ���E�/���v�牸{�x@z�D���R�U���t�$M9�{p-%��s#PK��P���\h���|��`i�m(��:C_�\p��܈ޫ���*�i��fX�l�ډ��{#�.�����{��3ψ	��|��2�{��<�>\�z�#�OB��8���g�r��Y��5�.r�%O}섡�<���'%)�\�Ēd#-������ՙ�`�)����cn?M��buJ�N?����!S���@�5k��^�ğ�g��8�F��T3��s�;=��V=7T���
�l���-ی�dH�������ਆ��ƫa�����;R�q5~�0�%�lD�"i��+<�|�.�M�;ŇA�J�!�:��>;uc��; (!ۖ_�V�c�����y���ȇ�^#�0>�\m��${�^�no(b֙��w�W�� n>�Z�>M�e��8۰�s��¹�N�ź/���~�#M�ގ���h�����k)� ����DЍ���}��T�MH�C������U ��+,�(�0�X}� E����"������o��"���㌖Ӭ߼%�!s]���G3���!r�
�#��-�O7�@#$^G�ڽ�9�O���Feu�'��dє��I����������%���,@->"�w+Z��6�Do̢27�I�,�
���H\�x,�D��-,3j���R��Oo�=.|�4��N��^i��F`��Ι����T�vo�
1O^�W8'V�%'s���`k#�!p�%�9�h�x#tT����TZ+Dŝ��ny�Z�[�5�W+��v��G����;��l����*��B5b�ZP��^4���6s�%�����R�z�������P_��	�}�T�X��w� ^���SUё�A��9��� 3.+#�4��^�	�L��!j�����X�U��T�����ќ�r�yh \P��-�ID8��[I����`�Y�xx��Dq�	�wÜ�U������U>V���4�	��.Q:}Int��,� ��c�&%C�.�����4b!�W�t,���b�M�3N��5^����(��5�4�=����/:���m�N7��͘k='�D�Ӷ+@��]YȬ5zv�q��JYʟ�n����N4�ڠcW@���� ؚv.�����d��͐:���]�U���n�a�;��<-CF��u<u�ԁ��|�PC�'Y��'�Wh�(�����j��#�����D��ML���:n:�O�9m���-Hz��#4+��e���p�q�1���r3�>��D�}�a^Y#�&����Q����4.�wMn��1�rU%aM�k��>~kR��BEf���S�_xM>ں��b�tD�l�W��d�����%/�	���&s*�����Y����I���{�<���־�U�`8.R��g��wsx���D��T�dv�jM;�O?fFy>Ө8�� ��Tr�r�\�>}��oI���NЙ&�sN�ױ�]Y.�P�L��,g�O&��O���h�RTYlJ�s����ͧ+83�o!vI��q4�?��vX~��:>��V��,T7�/�{%��О�z���g���!�˄��u4�P@�RJ]�\<�(�%�dMp�o��-�^4P��	j����.ã@�1%1Ӱ\��`�9��W_�f��K@o-x][&S, &�I/z�������2|o4�Dꤜ��Q�؄��L<���ո�y6��G�[{�J�f��qQ���9�*˻�H��u��-�qT���(C'�!17��Ul�Wf\�[�7��&� h]�q��-�vSEd���e[\����桱yE����V/�;�g�`�k��7Zt/��38щ��ca��|3?���C�,rO��{�����z���!�PV�;Q׭r�/��:�)H��%�����6�j�/��\�h�S��ƍ09V�n�vܙň쬢��&efL�-`U�&�s���0��В�.G$�����B��r`訁^㜟V���b4�&Wո� �{k�6�
B>��|'�oN����yؓ�||����i�K��+���e}W=�-��_�8�Cl��
�f��h������*[���@�k�YV<�Pa�䯾���74sC���Uk
}g�OC��X���<	A �{� �����$�@�3�8rxFYfh�#��M��Sv�5V�bBS[���"���L��"�]p����������0�U��B� 9��Q_����f���'H����J9��u6�UY�?o������ \_�/�B;4y�`�H��(࣪�>.�J���1���� =d�1a�����Ye(�'��e��خ�Y�|t�攱�g*�4=� ˞��=�B���V�e�lݱ��
d	5ơP� �^)жb?Jrne�N�0+�I��yn�{ؔWU�S����,������w�G����h^�埕s�my��W#ߺ0#ƫ���P�pBU��МܱT�r8�V���R7vԢ�K�)�����ɅƎD="vg i�#�L���x,�����]�Z�,�����߻�}��-�����K"���Z�Us��TVT)�н�_�����	��u
صKD���d��5�;��CMS�Qҏ�^@�D�4����
j�+��Uk��-�C�n��LUq�ӱ��MQ���v
.I+H��]�	<,���Ud�[�۸S?:v5%��[0*h�Kn~g,�5�$�g5��3-H��@�ha���?�]Xm�-ĞM�,>���^!����7S-V�[U�R�/7U�{Wz��U��`�����*XN;0'��t̛� =*!���b%n�b%Ea_�����6�.�ؑ��E�4���%��T��G�2m�V/#��7��lN�Z�h{��8��6%ƾPyv�P�i9w��eO���-�ﰫ��*TQ����X�	+��I�y��6LՁ�����~pY���2O�fya���e�s�
��K��p�|t�x͘u��^�/˟L>�;��}&H[y��j�����I�����}���P�|KX����z���P
�s�8c���q�`)	��\��w���@�7�r�+�YM&Ss���H�̢��b�:�*N�?Yf��A+��S�l����*�ZC2m0��:p5�Iaް	�v9)�,��I��&����!C����P	hmh����[B�%Q�Z�XpEf
\:��5� T���Z���c[����Eܝ�qX��]��W��lU3�LPS�9�E~�	�rBA���p~&���I�Xk�0�oV�Zş!"����1����s_���<�o��)2��'��2R������ć���~�9��E�O(vm?�]��8Q�W}�fhbEo�Sh~�Ы��QT��v���Ñ�@w�8�i`��l;U�a���3��9D>�݂�d��qc.&+�`�@b�(�&  Z��ڜfj����=���i��8?7(+AfdO��s$�7�R 9���e������l'��Ww�����.8h�T���ٍ����t!F����$@(���z�nD���	g��s�o	m<m\Qx�n�@�1b7�LI�?:��B੶�c�dv}d��ї\�>��
t�����@�mLZ״e�=�O��V���a�r���At�L^;9�⒋�gK.��K$�W���}��y���]I��H{͚�^������-傠� ]=Lr۫Rw�T��V��2�G"���d�� �mq��n�v2تi���٥]�u:+����L�1�񽕛�yL�	��p���z�d�����v�]�9�
���DX��@�E��T�YK�J�gk�'t��}Z�)�c�xdQ�� ��+,)!f��񮏘
({�=�Ƌz��;��6�Ob��إ���TEL�p�Ӷ�t��S������z���� ��+�=�����P2F0^��~ "����iA�e;��y\]{,�s�mg���8�/��r�O��ܲ$���x���	���\fJ(D���\�mj|Mh���έ[��h��(���](TQ9o��t���Y
�k��n�\�<ka���SE�+��		����ӽ��͉�E�p��<�����\k0O�n�q���E�J|'�n�����%�v���|�W{���� �b�F3̈Ĥ��'�R��G��wR��8�Lj��E�=�8l��qN���%T]*�_2:0���x=��I�j�V��H��ha����)�E[��i[@m^:��@�W�G�6/�pz2'��L�A������1���vҧ�R�����2�*��3����B�W�y�����5��a�̎Q��٭:dj����{�sc�.{I��$?=�<ʗ���ɫJ����2��"���~�Mఆ�=���L��w��1ʫT���c�^W���HI���� ���Ral#��f#g9S�:]���,�mIf}��M�8�Z��H9�3{���
J��Ek?�g�_��a��ӹMK^�QDw�^���X�rV�g����t�-@<�M�6���L� Q�@���[�-�[)��yZ)}�YEG�=�<���hH#ut�$[�6f1ȕNZ�]n�Gb��І<_�p�^��� ,���e�<Yaeٌ���rb�p���DE� �d�Ϲ�{��W�	��FKsV����
6��P��/�{���A�%m(�n�a�鑧2l�
	���v-�&���3uI{��]���������e���l��n�4,;�Q僗���8��"���
��	5�����h���;PGp�:G��c7��e��V|a�[���~�2�%��D�x������$��Z�q;���[mqJi�7p5����J�%�!j9۸���X��D�����O�`zP����w �B�8����@9kR0��rDe�#w3��p}E�����q#���W��A`*'|�p{��
ҳ�F҆$�[��d4�6��U| ~gS�.�����
��i�����d�e�����#��"ڽݶY@��7��Fz�ǙF�^ �CI��n�_��	3Gу:���O�َ7(BBvj�(�Ǆ�&8��HXK��0fV���7+!K�8o�1��Xn�0�D���6�- @��v�d|R����8�(�th�L���3*
��|l"E�Ҟ�eQs㮮�9}[���֫�Ԋ�K� �Ц�K�nTkȘqC�v�B3{ڛ��
�=�G�J�������E���v��z̲M��p&Eۭ4F���w�O���vo�z�"�Ir�N[���_�t�W[��3-�d���I��-c�rtS(yh��6ĭ��6ɇ�uJ�恤�O�xxDH���+S��np��|�l��p�3������~�l�6b���/�Q�W�?!�'�2`A�ً��-~]�������O_����	���T���Zt����5��=��L�&���W�-]�����j��C�G�1##������q��؛8�u��P�q����钱����w�t���2�K�8����n����-�tG���ɞdH�F��;��Kև��$����i��J{�r�*������Ҹ��;K��&�ꏵDZ����!����En�[�3!b�m@���.f��M����Ԫ�,����{a�/���E�`�?}q綐W��H-AJ5{"2��7�9��m0�v����	014:��˷��Ĥ+�;��\?ZXi@_NRZׇQ<�c���h~ ���?�*�F��CS�}���Z�gT
&`h����'�I��gӥ���h�*f f�&_�#�p�w-���F��i�շ�i�����Y�Ŝe��)��{�~)0�޼+?��m_�6�t�n�6'Ƣ���\P�b6y%i���_��i���̢�%�� }�0I�b���P1����BFE+==�A�^��,C�:�ظ�
Ƈ�)���'m�7�*x�h�9�Y!S�a�����c�|��yCW����2����Ǯ��+>��hў+^N�B� ŵ���O�`���a�8�a���Jx��Zu�L���&������o�}T�vފ�gGD�yT�:�-F+]�D	����[y��>I��cH��DR�U�)J�Oi��T4��2�u_�v2��;�Hi�
I]����0��=�\ ���*+��r���X�Yg
W�#Ε}Ԕ��H^̾�g}~@4O�9���d�n��G�^ ���
�$�mk�d�ޓC�l�>93`U7K��5�?�9cc��}�X���siU��G����Sn�ՌEk��q���M,�7��*�+\$3{�"�Q�v�6+n%�7���s�#�jf��T�qU��H��z۱�>�=w:��:+��S� ��-���77X��LΑ�Y��c�NA@�B��B�!עơ[��zA�"{nV���j�g@!7t��F>�1zYro�f;���#���@�q֩�n`��i�Q*�,6��Χ�W��RTɃ��.�%�Ǎf���yV��2�0d0�a���e�)AEEx1�KT�o��g��66�g��M�شx8W�X������;�6��c!je�-Ó2��b��Ν��R��-z������,������/�JM`:%�4��<`?=or��3��2�͈�a�s'DbLt��凈׷�hl�5|����G�����-����9M��>x�P��q��"�؅'�Y~ f�o��0)��&�d���b �c���o7�5��VM&>&��p5�]��M��η�v3��g���ͻ�;��gcF�)�Q�wk��t)���q��\�2-��@�H�3[��Kp�M<w�/G�o頟}0�CY�x��b����)}�ng�}�sBhB��7՜�g��D���l\m����g�z ?i+DK[�aJp�##��	4��[ÌW���N�u�搓&�=|��g��zG�=wx���ed�P��9U���0���(�ޙ6p�޸,�c�=s���a�	��3^��FD�ZG��(�0{)���`�0��Y��W�ndQ�@��.��5��r[ljVf��9���?-���P��}�N\����ٰ��l��b�o�	��﮽>�zvP�>~E���ʄ�T�9ޚ�~�!�8P$��Iwo�O�mIƨ�+��Y2�ГC��X���HࢯU���`�m����CM���Z�W�y�$�c���e�<�������_���Ñ�P枙ƩpBtu`�i��A��X}�@���	�����n�s����4$R�������Qj�|2F,��w{�=oA�U6��h=D�j�E4%��;�� ���:�{�S/dM�3�4��<���۝�I�����Q��NȰ�"�pIRxE6�0ۺH��Q�FRKʛ��U�q�%ϓA���K���~�z�s�ؕ����������В��*�6�kf{��r�&�2�T�̛i��^��.��^kS�8�JE�!t$�r��A��`�)5bC����}ױ�gW�B�*�8�!�[�#oṹ##q��M4j�=�m�?��9jVX-f�]9�ܕ�����%+! �)�Jj�� ���GDٴx$��ZQ2�;�ao�N1b6��X��a�~O	�����_9��Z�&9���2�%���p�eQ���xԏ��Î ϶��K�|�����@��l�Mϧ̴v�/���Fz_Cz�����|�^U��w��}��Lz�g��H�~���O�3� �������V��@�*,Sj��t;S۶��7���T����u�Y���'��"ݤ,� ���\��?��իC��m�2�A�>�C
���c���q��Q3t�i�CGWL��+���&���V()�Z�7:� #���+G����C����8��&ok���fqy��JP{=v�P��:XCVХd�OJ���6=)[g}�C��d#D{Q�J�M:����f0�����=���kޢL.V@�c�t�Sy/M�^���E]4�� �q��^����p�����h�\uP&[��v+��z�����y)��p	���V����F�rO2*K�h?��2�T�G�M�|{1�-�O�MO����1O�G��"�G'�~KM���	V�\�V.�/��$�U~�k���O5_)��c;���1g+b;XW�p�~&�Q�Ӂ������1�fUg���Hs����a�橲"�24�BȊD���w�!7x�|�AȦi�[b-�:U��@ɋY���xqlIn�vh��L`�k�� �w��9������E���d��j���;���"b`��٢h����هY �Ld.�B��)a=LE���c�z�{j�[�����:T� ���[5�xW^���T1Ұצ@�1�&/��?�]�q�k�2Nxql}�K���͝m�5F�EN�˽h���&�P�hߛzKii	���uq���r�+�\��=�Y�Q9���(�6������®����l?f�	<�"4�T��3͜P����g�Q�|�e�e9Зa;@.�BQ�T��� M�(�t04+�,t^m��d��C�b|��tzS+Ab���s��1�����GO�[�S��lfq�<ӗ������SE"�D��_��m�����Q��Y��-�R�����3g����]�`S�f�h���d�o�A��q<̾N�]]�>NI
�.�y�$ب����\��E�l�JG�[zԨX2R��h҂{���7'Q�h��?�NjCc�Y4 �p�{=�{?�C^B�c�IqX�BdI�X$2��1k��,��]޻���=�/��E�Z�,�mO�
��Of����&���3
vQ��>X���y��f����:�^޷u��|Y<NA���?I�ҳ�y�;goO�h��uQ&��Ļ�0a\~�ҍ�>('��{;^X�&�e��%��!*�6����0"�2�e�3�T
zÅ�_"�`r �: ��{��Y����Ӟ�F����/��Q���ю|OJ�ʽ�G�õȆ����0Lik���ǜ�c�za���Iv����&��!![4�A �ИS��iSw�M�*P�O�/*�%V�V�:�Q/OF�c�s��]��<���[��Yi7�����f3����%w��ȓ�s�VL�oJ��
�	�"�}�%$��?"����!�z���(�+�B�h�7����
�~6_�$,�����Q��A_�;� �dw�?��&�_���E�Fp��s���a�ߧ��:�r�h�[(�=7kg���D��>��ˁe�P�(@� D�p�	k�%CPx;���^��F�R�Ku��w꬧L����v��I����Ho�#o�V�*隡�z$���A,��πBi��	�����"HQ��<���]������֍�::y]�֬��(bzj��Xˑ�!����/a�)�az=P�`��:�S$�&��Y�M���>�=Hٱ�Ҧ��9��ٹ�?Ў6pEyH��Xhf��>�]�$�����/E�f�@����&���]A�
�K��d�If��	@s"��7z�.yW�r>I_�j���+Ud&|�GO8�HA�yV�*��@���7��V�i����T�������1c��*,���Kby��a5�t�.Os�<:�~m���C��?�d~��=KDo�WB�sV��a^�������a�1R�����v:#��9�u���b��DV�d���4S�=2$�&?��u~�N�q��m����)�ĉ)>��A��tcI��&]�ӧ�]䅾XN3�hF8)�P�dX-�`�}v��i�ɿ�Wjs^4�9 �}�s���"	�%B�ֺ����"����
ԫ����U�wR�:�����(��[al�i9g��EЛ3��%��>���Xc�]�J̭G �_u��ϑ�>#ĀXq�~���F㝵�W�����	4������O�$?��$A�(��Y�*�P4�
���푾k�{cK|������D,ts>|�d��e�Ȃ�z��^�_�28#��|z��.\Wy8�oa�&[M����W�Ƿ����dV�:0m��vΐ�cZF٫:ാ�X$#,F�������
:�ҞJ	N� g�ũ-��P'���wߗ���N��*�7�Ͷk^~H��)�Qs�~�Jb�}��⪟=?�6ī��Wrզ���j�G�Whml�l�1*�����ؚ��n�����n�iơe�D��>��x܇u���RRm
c�V��G�>��!7��*)��sx�_>tN\C��xre���?���*+���r=��[]϶J��1�!�27m�]h8ټ�F0E��mp�����ꇢ��u�����w�RXZ9VfOJ��h�a!�CJ�5�o����g�b5)&�>d����S�U�ܒ����r�]\P �ܓK���3�?���
��M��}�3�����"�N��*�Vنf	.�3fZ�ι���G) �=E�w}�aM��l8�!��!�Jl��f�2q��(HVj�	�4��f �M�eM'�����X��P��G���y<ƃ�V�b�NFm�E.� ��O�![Qى+|���p��G�?�m�/��|�	�/Ԥ*���Ӧ`:\�A����� ��=�5�h�A ��O��}��i�@Dمx����88��#vȔ�g��]U:�R�`؈M�$���xx�O��\�}�V�`G`� �u�(��y�6���H��^�A�B�F�U���u����x���V�s��7�]�$�ɤW���UH]��:���U��+�Za�F-�(��t���
L�F��4�Ǣ_s�J����M�l~I�s�)������3����iHу���o�"�瀺u�a��vɦ��VP[�ڮI��pJa5����
�Ҹ��f�ORB��
�M��H�vp�	f���VYS;��R�>����vh>����a0���-�ͫ�,هp�,��mى�����O۽�3ت�)"{��d���|OHi6�����eX��$t��Ǡȋ��H�c��g����%���-(��U~3���*�F(5��V<.U��>k�8^Ee�.ۣs�����<���u＄�Z=jRFr���9Og\A�9\O����(Ha�O���8�������}*��'��
 �@���oHj|�:�6�?�WI/Œ�n+����s�5�]p����<� �\{�z��ԮlØ%ś����?�E�H@m2�y���p��)�[n����#��A��m����"��h*%��}�]?!�U\Ij���������LYNw��h~��g)>��^�O.�ǂɋ�+޻����,��֔^�������Qh�	�.٘Of��6`��?�1>�գ6V���YN2�&��ۥÆu_s�K8�c,��"�eܜ�+��*`H��� ��1D�
r��dWdZ6=��ap�Q}b��ad��c��S8x�)�*e	�6��H�Ϲ恻ݪra�|CL^=��s]��f�*��;��l��a�{���Ʀ�:c.)¹���,���
_2^B�^�u5��HP ^v�����1�w9�g�C��kF�7�
liWA��[�~�ռ��
���޲u�C�5C]a;�����Ø����eq����;�"�W��ͫ��Pz��qbP1󫑿Bi���a�����g_���2Vb��E��)p������(F�\k�oW��1�X�P���ޥ�����@bf��6`0\�����5��}nN��x#�4��.~P�?�o��q(��9�H��j)���n��|_��w¥�?�d�O2NL
墊�i9���ݾ.~�
8awR�e��"�,�%Wu�Y�oA;��ԊC���<@�.h�D���r�"?�-)�H�>��ȉ�P�YU��3�D���\x1��(�tPƶ�as�f�⤦� ��x�{4�ˏ�ǁMtI��T���{ŉ[ �}����K��mf �CT|ԧ�����PpU��=�g��K{��AʦJ 0"��i�dn� 4*�_W�ji�큟�v�x/.�P���(tDM�x���&�
s3�J�������n�?[�R7D��2
�,S@��v�{�Ӑ��;4�3Tv�Σ�Ͱ��ƛ�܅ղ�kbr�{��*%R�����7	>��
�a��h��eԾ^����,���n�K�����
�1�v��|hf����Pd�͉��ACZ�)vM�Ю����r^e�E~m|�Tn��⩆�se���) ��ֿ������>mj1�����Ms���Z���p�����p?Q�_��}ma�f�U�F���o��ܽg{����qܝ)��v�#!�8_w��&�+��a�_,�O�F�,��/?����Ƣt�S9��:G�7M�$��obX���+ԋ��_,���l�cp�Z���9&�:}y��/d�-�t�T7c{��z�/]"�6ݸ�I�{������<w�k(��&xK�RQHuJC�F�ﬠ��AuIK�T}B��QV��c*��p���\�G�$�?�VL�d�H���X\����̘��Rts�ȓ*�x���R������SJ��E����Gq�P,]�0��Xq��8;������%Rt�UM�_����"��]�)5-v�`�0|�,@�
U���q\��{�]HK�ZG��8e��o�r�Z�2ྚ��[L�LH���!-c�g����c�̾�֤���������^���ݟ4�����\���:��9е�����{����w�?�朗S�`�L�ed�W�aք�;�ܬ8�'{L��!���I
��`8���\*��j� 53��>TIVX_S�m����]mj�$z%J��f�x&��S��G�%����������k�Y+��f>�|� d��k�ÏŲ�4�Ȥ�
�.���������.��0<��1�Ix�"w�o��~&����7�C~Xa�=}4k�yԶ�v��S� ���|q/�Ӑ��;����Г/.N���XP
?5����s^f\�#3m�gc���)m_iF-��7������9>x�X
��2n�ǩC_�U�f]�A��8Z������H��i�VjO��E��ͫ&N����������}��zj��k>E�J��bg�y�W��5fb�[�?_��^�P��U)��}����_�ѶF_a���`x��ޜ�'���!���Wd���VCL܉wܪ*��\����&`xoRr��/���5�e���R�_e� lj��F�<���j!��_��V�.>{���������D���ʱb���r���zTP�^agt����~׮���QS�_�j���W�܃�7O��e�6VmE"kD�ׅ���Z���c +0�>��w��R��[���_e u�lp���ٳ�6�u������f�7DDE����J������|t�c�Gc���Z%"t,n6�b�øu*�*��X��DMfi[�����S_�Q�[P�Jz����B��D��T`����oX7�	�k�2�T�.#��U�rQ2�W����!z���v���Ҏwu����q\�U��l�
��KX́�(��A~d�����+�ڋ�VB���b;.^m�UY�v�F2�7soR�@幛h�s�X��+��rboc4���d#���'�)Ò�oɃRǻB���z
j=�X`'�N���N��`R��F�Y��~��M���5ZG�|���(�Ҙ�yz�X�����S&�b����!��������D,���onLcB6R?�'r��B�o��������ܐj&Y&r���7�j�u� ��a�D��A�&��X�d�nr�M��I����<d���9lm;��	l���'�*����#����(Ȁ�A���8
��bZ�rlg��
1�>vɇ��f�Û�^�{��ɦ�X"��]�&\ڂ�b!6>@�Ժ�j���/�f�!�JHH��XpmW��w���������Asb��KE����Qu+������	�t$����?����K�``���ao��j��d��}�c�nu��[|�o�������J��^�`������`(~�*Q�m��������h�h{��� ��y$�דz��c�(��MU�����1t��f��l)]�C���s|z�re,�W��=b��j�(��$̫<��o����O�j�m����hJI�z-���W�j��+TgPW�9� $_[i��P�C�̪-��	zI�;u�����A,��H�<8�d��3[Htr�b�{]�>�[��A���/�8�g'����T#������`AU����Κė��l+3�ۄi>��I���})67;8��<����+�u�����q� ����IF��Y��!�N�b�x���آ��Lۑ�䝘� m�1n\vz�s��#58��U�� �=S�T�"~�!�Y��\I�B;�b�y{½�~@�D�[�ևEw:�Y|Q���^��Y���~.������Pm��k��9�D�Q���wTȉ;@�H�NX+޺?U1��g�H�1�۱���e�|����y��G.��^5,kXjӵJ"�����+R/�����V�P�޾�ǜ� �E@�qV��Z��oh���G���y ��X{{��X�%�6B�;��r��ð��l���M��O��?�K�uq�L����?��~,�3��;�A�Ix�ϓ�X�#��Ô��?*�Jt�ÿ��c92��U��C���C4���W�8g�̕z%S����p�ލ�Í(c��VU�8�#0��9g����[�2���<?
�J!�Y����	����}��3<�z�vK��rB��3�1w�7dwJ�	�K�rj����9������V�u��e�7����y���JT�ucԉ�.�g=p��ѧ�VgAb6����`J���W`6��`3_���z�V-�#��f.�y$��*�&]��g�w'_��������1�a3��5�������Ӄ�2�]��#�d5'����'�@�^e�G���k��vi�k�-�u������%�wyuPA�M����#�	7Ȍ�����2�č_R�*[M�AZ42���Z�ȟ82�+`� e���8����|/ ���I;3����μ�����xڴ��.���+D/��H�A�5��ଊ�x��硋Z[(	t�(�x&�<(�	
uzY�7����O���������R��6[�v审4������o�V�ݟ��E �f\'`�5P����j����I��ܺV�~��:��a�BS�_��	u��gb(�Sc�60W��̏�ό�	��Z�4�:=o�/5���\&��P����v�;A��+��,wB�^�=��5.x*e��Gb��)��e X+�L�_L���9��@�v��M%��5[�v���Q6	��u�Df��oUW�_�"�ӑ�*�̫$O%2�m�l��^h���̤u<M�$T��� ��qԯ��a�h��������qv#���h����N�)�i�	�dp����`&�o/.p���P�8_��N��H ��Y	�Y��ѭG��������cx\^"I��2������zy�t��3ت��V�v��'�@� 
�ɛ��ǆ�tDH�͔�`��A`���|� hջ�C^W���O�"�!+u��M+�hZ(}�s}�H2�ΊdΝF5�W>��r�s�i�W�k^4����_�p��e����w���\���5SX|	F���OR&N���w/��n1�@9O�oj'��H>�"#�9e,�2��t���x�I(��i�-�^�����|����/����e�iR;y�]Q�ZF���U�T��eM��*3:�S}�pvT@C?�F�JBI���^�G�ݺ�b��l� ��`F+{�q'�@!Uڬ�!��UXB/T#;�_�0��M����'�m��)%��V1��M;R�ѣ���6��[-��J��,��x8ăh�X=���ݳ�L��*Riܖ LP��lyUuJ���S�����_}�Z�*����4g,	�{=U�֗��~��.�����7ɒɄ�%���&�?t�v�=Y�6x�DY���O�nݒ6Ţ�0Cw�V�Gd�-I��\�a��޷�\�������<$y������"�:�,���np�Nwu:�bpi�%Յ�eg����{�G�}�3R����!������J��lҜ��]��s����9��?�k�H���T4qB��o#yQ)ёr�`�!rӠ��B�m#��N������'ژ�C��!*\�����u�6>]�'�Ub����R� I� 4ʈ
 �\yѽ��=2ʀ�(��y�6� �x��� �/8�:�~��j���mPk�ǘ��,��SsT�^���-iU}A��=���/�;�c�?o$�{c~h�������w�(����(7<]!}(�[�t��Mz��C�)֮�M��> ��!�ȯ����!���'OŁF�:��R���0\�zE�%�7��CG �׃f�O��P��݀��~��5�zcM��H+O ƻöM� �3A�#�X�p�p�U��;q��3V�]أ[�esB��b
h�pF����ܑN�֧%Oޯ{/���x����� \��q��� ;߈xi
���>��iʽ��ƌ��J��CU«1w��ܣ��w���$r;M��(�0�i����$�x�e�=�H]��;�d��j01��F{�*ٿ���X��.�L�]H1jή�p���"l�'"�p"ب�*��(I�U�����g��ΰ���_�̈��p�n|=OR�I��%��rq�t��m:+�¸��k5?͖;��`4BH�{\����.�������!�#��s�I�0Q�(��`���d�C�0I��c�]���?A0�dF�s�FR�v*Lt��L�w�=��ښ����%���	#�ByA�gLZ�ǉ�e�W��x8�^&��J����?�#*�8�`Mp���ny��(�Aڍ�oڽ�}�C�U�4��^<�?����xP�ʐ���Q���0����s��e�g�GG�iXP������2��_>�����(��`�B@"��*V52Z�2�nbUE.�;n�o{D�'ԁƪ�>�E�;d����^ė39�1`�g������
���%�y��ty'r[K��-�1 G�t`��M�W����tMՖ� ӑ�8	�&Ό��D��.3]�"��+γp�.@电����s�O[
`��\�z�y(�7��Huڇ8�+Y�,��C���4��I����`}�;����Q�u��3��
��T2�k~w^��~�BJ�<�S������@@v/Le��k�W��1pt����L=�r�yDjf�ŭ�/�Bkχ&8n�BR�8 �s��L�����J��ŭ�Sd[�U�z�(�]�� R�N-�oK:�p��Ec�Wԣ�Q 冧�=a��,�eM=�tF�
ʔA�H��7f�����ľ��
��oF���֡j�<I�
2m�ν��b�W#z��ˮ$:�>S�� �ӹ� �Y �7)�Ǘܩ�[��s)D?B?�����`���&C���ĝdw���Q}�}T4/���Fq���5e氄,�L�p�_%ZjB���zx}�lzL3H7��q%Ɋ�,x����O�ص��`���w�R�Y�&P��*�nv�K��Y��w��G��~�E �f3�5�����]w�J�����i��3��i����0h�
�L��@�K�^�)V��n�^�4�R^s���rC�U-X	m�\�,�,c�#˼`�E�����"���W
Zt%G�$�_�M�����C���y��z)��n�k�-�_�T���S*B��j>�}	 �R�pM�F��.�*��2�ymo�6�Lyq~��2�?�o	0��m�cg�x�D���WVW1̾�u�*�^-lAd����#d�B��?�7=����衭����>��� ���Y۔�I��m�9�0MA���$�ŝ��b�s��v)7e�~	�"e����b�ĩpaH�Z���^@f\c����L��N���l�0sOQ�y�u`�8؛�nN�}0��8nZhB�Q3&g�� θ:Zj�(&�v���^FS�,h_^z��W#r//�^(��H�%�g��S�c�
?K>*J �
����+Ň(�Lr��	}jOҤ
G�I�W������@���V�E��5��^�ro�8�����M ��݆�D��y�Li�!��{�>������uqiY{-�>u^JŃ����فIڇ#�R݈龄�ÿ?��a`�1��I�(5~u�mŊP���輝����4k��7�!8�uMp0�/
�lq�)R9�L�4䙎�������GM%A��A��	@�E��6���%���S�e/x#+w�!7�+�6�r��k�i �f�h`V�8���{mQ^��2�����VL�pq-HS��J���߲i�A����"��o��	��D���UӨ��z�Yx���f����>���,F76i�)��{�o�Y�$���x��l6��K$��u�Φ����k8Lb��~4�IG_gj�` �X�0�b���'���h]����M{������g�K�_mo���,a�6o'�U�m��D��5�����1Y���g9L�Sc'�̣���(�dV�������[�9"?%�\��D��i�ؙ�����mD	� <SLr%�SޖoO����}HF"�38���!sv��BpO��*4h��T�����NK�������dg�	�ƾX��.%�s�`�?R�"�Y� ?�ʲ,�A(Ln�����Qmۺ:��*5��]�V�/��'R4��LB�ܧE���|���G�^,����{���i�]������Lv+`![Wp�f9@M�1�
!�Nw:�q����UQ1L�����ٔ�}i�?����}D�GY�ݞ<L�COA (�A�O��99m���ɺW�&��Y���>�f[ӥ��:x�ω[�xA��yp��-��Ϫ�!�u�u��iF��tA��n�2{;`�U��*�
����$���jOtA#���ddwQ!�7��/���+�dڋ�B�0lV�����6z~@��u`mJT�4�%��1�Y��Oa'刀�{�!��O���$V8�J�E��	$Dxb�Y�^H��9*U�D7����TM��no�v��J�`O�.͖���s�����Ŷ��*z�7
�<�#mM�5������T<
t�%�~��6��v�2Q<������"��-W-�L���h�骲¤,R�T�Z���K�ww?2�w�p�7J��h̹}��}O��7?�&,\�tq���f�ϴ_f@��㶡�H��j7��v G��T�/�\�Wo�sH#�{]@�d��0��uR���`��M�}�ˤ~�h��h2k��Y����6L�Q�f@�3l��ɸ'd�f� T�G3���=p���=����t�7���T�P3O�V����X��Cs�Q�1��X�6����|�'�7_��(��MJ_�[��Q�g-H �1��PH`Op��t��=�Xc����QP���z�Ѓ�]k�����R�\��/�Z��8d<WN���˝'���R�]���N�V¹}yS����B��B��צ�����wi׹F�\�y��'�|��D��JI%��a�0cY���� w�p�}��Q���62�y.���L:~(%�ڕ� �P�X���y��X9���;	bO���)��viZr���x]�u��,$�|�>�I<�hMq~���g��J�e��z�)����){��k<��ݪ��� :?������'�7�0��7)VM�ڈhV�H;��!����*�g�譍��@��k0Z\�9�]dX<�g���ĤY�|�y�<\�&l�ѥ�X���M!���ȗN,�M���A�&�z�CfԌ���_�#���Q2Mi�����w2�o��?}Щ��lG4� �A�K=������nn���y�^��/RqA�����C1��Q���5u��賉o�Caݩ�{Q��x�����S>&$��[Ö~��m�r.8˸���)�Sk�!�x$�Q.�e�cf�\���S�_w��V���ᄀD�9᫺
0�PG���TlHyҨ"C��Q�2O��������g��$&��ApO���W��[�|6���d�s��}5�2i�┐�f�7�<�aN��͌��+P�-4��ݲʁW��)I�6���׽B�U}�3sα��{2�Q�5~��Έ�>U�k�r��2��T��Ƃkߧ~�Z5~������ ��G ����=
���
|�.��ؠ����g���R����;&-�gK��5K��m��%��a. H1�R�LU��{� xyGk�x�	����.�����^�,�K�Ng�7
��ү�1Ftx��m���}���3�x�@��{$�e�/q"vH�I���ÿ�Va�pE�a*ϖ�X�Or:N*�we腰j�r�@�k���,�b{���N8�;��W��_A9^��b���O��kav�kEy����D|MBw�����Y<��A��A�����''��"�����W���� ��7 X/��5�t0�LW��E؞�A�;��P,m`�e��;�-����c�R �("�	~��S�k�K�I,1{5�t��� �_�,���=�#*��#�ǯС�?%��K*��jn��������G>�H������v1=�:D9)
���'F����V#8ʘ]��[���<	IR���n�g,R{��R�T���V&ϥL�vѦE��X׫1&Վ-6vZ�?T�{B��_�n\�����^C �G�v�o��ꭄ �����PtL��.�R���ْ\�k�GC�d�7�@{�	�������Y;07���w�c,���O��D�I��ؒg9*��)��ƾ}~���?�E�Cڮ����阴#H�BSCA�n�r��$B���9$�x�C���xVmg��}'n��G�O�L����;?��jN4?��Nc�p�8�oy�oMg�S���{�0|R�6���������W�!` G�T��	���d�[+c�]B��l�;D����B�Z4f�Q�x�9h��=�Ⱥ��)q��+vX���m�#�,Q����%O-���`��Y��̥K�x�r��팉�:/!9*(2�v$�W��:L�ё�n���kw�Gl,�[F����K��

U���&ゴ7�ddqX�D�AD4߲	��+�#9J�z�3�����Ad�X����I�di�Wg�~�����"l��@"���Z�?}�,T�&T�+6\���b�	&f�{C�n�ib��倌������e:`Wm�T��p�gp5}U�Rٶv�wB����$k���DF�}:�(q�J9'+����*b�td♴72q������y���r��S��A�+_�4�߇$+w���8aH�����z��$�y\v-�����!w�6�(��@�3������c%�#�ʃ|7��s���U�'��U!�"�蓡�4^�������4�ǿ�Q��?��5�@җ>j�ha�ES���.�"Y-�/��j�"d�Y/�Mi_��.���i�X�g%9�$$b-!(>���I~��4�nxS�������l�#-���_K;Z�������$��L��l�s�ym"�z������F�>�_|�cHև�m�çj���gĦ��k�V�K�&�{��ݴh��2�S�|��K@�ë��ת��s�J`�V�x�?�wv���Z�,��FfR�cmeZ_���|�f�a:���h\ڝ�)�Z�!YG�ca�A.P�)��~
U������2T։�U!���ɓ�b2+�n+C�~Uj��m ������i����l`b�6Ɵ�U?�<hPv6��`���/i��Ή_H����"�o���{"�^!��P��~SV\W_�#��;�"�BeL�A�q/�o�v-w��/Ls	x:L;��h�f7�4ޒH.��ln�T|m�]lr���1NW ���C�0�@t�s3rE��4��!e�}+�a�~Z	����L��� ���-�W�ͭ24�e<��l�2��6��p��ł�d}6E3c�K:�S�����U��3���s��E,e
�S�r�hP$�s�U>2���� �ƺL] �/?�$ �{��RF���\����G!�� �fuq~k��~�ݤ?�u��Ӝ�	l[h*�����Ma���4Qv1�uVC���̴M<�;%`⋎>h/��h�?!q�@��E&O!��׺��H>f�D����Κ*(�bmW5 ���	Ɖ��z
�\������X
��Iwv�k1��q������6	�LΖ:���[�/kP�*��$4=$�[/����j��Z��ډ4��VZ��S$Z���U#�dE����$���FB@�/�8k0����K��#�ô��X3�K�Ǡ����w��X�����4����6&�	�֊5v��t.�m��Ư�MU_���e�E��V&��ocB���ȶ T��s�#b�7���%�.u���<>��&������`�����#9�����wg[B3-К�?hڥ��O藃,h�a�X5��ʈ�P�P"7Ս,�qܦ��W@z���.!]�	��0	a�8��t�vxπ��v�j�2����m�t�) ����)�(Q^cz?<�ɧ�{.�£<mӡ�f�tkeF�s�	g�2 G�;�ܺh(��_rQ�M��}f�/1�3�lR�G�ؗ�Q7R�3�H/�z��MW�y��Ê�mQ��t���[�<��eŇ/��}fhǰ)e7K�R��wv�|ANC�+	�Ʈ3��]��K�!)f<��,V|����z -Dy��1�&Z�/G�I�AJJrԯ��O�
�7�������ײ
_���l�C(M)��~���s	jv���y�BY�9!0|��
q���3����"9ݺ�q�-�
8� �#k�m'+0�AJ��Sz)��������8�!o���H�h�~^���S*��yO���3{�
y�(��:O>7.)��f�^C�Wjќ�Ų����o��ȦtH�@6Z@]�|�	����d�R?�d�&����a�ED����O�|��$ x8��-���nVR$�
�Q�2c��'���9���^ǧ�Ř�Q�D�,�_����m�k��������'��tL}7$ێ�NB�!S���Ȋ� �K��W�	B������M��a��F#9��=�P�j��3L6�_2ods��瓤1z�Cv`̧U�t��n۵pM3=^�v�Xؠ>��xmؽe��)�3�����S���HX$K��o��n$Er����Ma%���a�[��j%������Ȇ���N/')��Ć��g��~�Js��_��sxY�h�ĵR_��v	q4�ÔX��Z�O�xMK6���,�'0�K> �ucz���Ę��=��!^o�:���)�{,xB��^���U�D��1M��6�6�E�/}�̦~I���zm�M������	�1u����&��F�x��Z�*�8�#���j�Мr��&��\O$�H�%�<�G��>-��u��R|��5��'+6~L>���� �gQY���j��Qf���oGs'�/�@![�\,�^R�c,�ԓ�6
>�:3s���zH��W��E�ǌgW �"�T�
�I�g31���QT����7����g_��i�7a��bk�������樻l_��2�x��F�uч+�����A����XT���5Ā�I��`�Ltm#I,�6ܕo�|�r	��m�%��~����2
�NI�fS�����"<O�#m���nT%��#l(#'6�n&0��2�Z1�[�i�]���g�1�`R���kd���
�qʚY�����[��t|6_�}�2I�]͎��T-� ��0�zY3h��;��n�2�Q����x��p�`��������l��m��&5������r)Z���j��RVyٌ����j���N�|�?�RJ�A��\�8�Wh��c��E�$.��YKI�IϻiJr@ѵ��FA���)�z8�������U2p�c���-[Ԣ007�;�{��V��&s�_R{{20Xc�{Fv�yl߽*f6,�ˁlUD�ڦդ�HˉF��N�17_;=���*�.lj6T=����O,A���,�����0r\��ny�����NZw�(��qn$nj��]������Ev	g0z|J�����{�El��SN��ő��}※�#�nm�E�	�l�s-�忹��0�{J�+�P�B-�0�� p�۔:�V����>j�D�^j�#W	[��dlY�ͣis�g�uF���U���͙����K��"����b� ���%��$=�gk���4h����C������:yn�*/v��H`�������C��6)W� )PlP����a�����X͉놕)r��2KmCi��rE��4�>��[��VP�୧P��Q�e.���>TI���\]9��kHj�k
1x�3,�zP�I[�.�v��
�7���-�d��N���Y���icz���_lu�)��X����#4�ѷ��T0&���U����`�Ub>G-��-���%��N�u3��τ�3��V���mэ%�o[������F>
�V%�Vdq�l?\�,l����i��^#��P��L�#cG�ٿ���1[�/�	9�����x�tc��e�	�:8u�b��dH�E� [ ��\o�wm���mȐ���90�@׊S{4t�IߎΑq��|��xJ��uTt,�#�+׊v�@�*��x��9g�5�<Z��/���kFhv����X�`��OD�ǃ��y�����^o�Oh'�tgG�eƁϽ�b���B6.�L{eOh<�>��	C鰤�����D���xO�7��hX]�"�U_M9n��G�;��6D 1�\���0�␕t�N���d����H�1�==i�;��i�m�E���eaC��?fbL���ߏ���`Š��9�Ԩ����!u$͌$��fÉ:D����uK;*r}�m�kIh${c�
X���ӸR��$9cW�=p���9��S�8�I��%�c�ϑ���Zʪv�[��[F��e���T�T����Et����R�7M�CYQ�(}��%��~�ޡF�@Zf�yb�j���D�y�N� �-���۲��^i�P�7�'�W!���ӧ�sԣc���#m:�HĆ��X�N�F�D;B�̓/���Wx�� |���~��#�Q"�X��2:���1�n��_ow;�e�_���{q7YU�c~��Ӄ�@T9�7ڒ�A�!2.���`�;�S�#ݟ:�$Рjb9��ww��e�u�C�
6���1a	��60��S��i�w��i٘���Y�9]�Ŧ@Fp���מeL@�GhM�*�TU ��Y�I���*wB�:�����b)�\��H��:�zrq��~����]������n�<vk	7��C�x��k!LS;U��GA�6�*ºhE�S�R�AG�:i*����=.�6I.��yt�J��O;h�� �R��'�i����0�D�G-�%øHU�!/�	 �ܘd֋��RD�C��ơ�7�&sh�� v23�J����n>%	E�/�[�#aexz%�Fz�1.��+��#v���pܾ��dxy�WT���
��O1���.����-�ZL�Z^Ծ���͙Z��S��_�i��7�q>�Xx��M���?� �	K��_�ʎnQVr�3,!}V��{{(�����H�U�y�����j���U�y߶_�>�u�{�ѥg7
���[&���S�쁳��RZc�:h�>����0(FI@�!�M.�4;�Q0	f�\��V�<�� Q�K$.2��.����(qC�}<je�<�f3B���}A�'t�˳`���J¢�)ټ��f���c�Y��εك�*�&}�7YT��n�kDˏ�1�Ǔ:�|�������%ݜ��].���4+ �mi���q�y$`�&�8ŵ��s��H�,gF����v[5G�T��q(-0}d=�S���s�.�d��B)��:����p�Ϧw�n�I+ kea�lj��E�K\. 1	�u�8K=�L��nY��;��V|�umF-)�nY�	����o��3�y��X蕶+]�^9ERu}�XM;�~�����Ma}���J��X��.=\��;�zl�H@���ɛ��3���ew���M�)� �͍G�����jng�g�-b߯VJ�'�㯥�=� �P��@��h�e��t+R���Ј�(�.�,��5�|���E���za{��ۛ���pޡ�L��þsSˆh�g�&6f�N��O�K%��l��b�)ӷ:c��~�ȥ�}���#$�ǣ�7޺��<k=ãcA[?��%W�
A�I�E���]
�* ��� ���&>0��8$>�J�H|$"i�:�~V5��-CU:�刼�t���Zs*Za�4��]l2�~:�#ƇfsYNE�5k*����<<�y!�b���w�$5 ݐ|�Մ�2nǔh��o��:B�Bس%�����O&�lc�W;'��s;��:�KI[�_�%��Ӟu�6��L^ZJ�{8uW�@�Y����+h|�!�@��V?�����!��B�@J�=\�6�	��D%š=`{k�%�,�u�'ݣ~ �ʉ?�����C���O�����C�n��enǶ�C����_L���zn̴T�kx�C*�0)�?|p�U2�ޝYG�ύ�jgAW��ë܍�r����lg[�#
.�N�L�excԌ
���1ȢY��"&�@����S��w�<z@��E�A^^�\y�V�~!�T��27iۏ���˲.6��70�s�5��@�&*8�/�D���Yݷ��K@���T�<���#�N[�.���a�9�C�h?����+l1 ���N��Eh�_�}粶�O���!zNsw$L?�~='��Qj~qi'�v��}������Ԭ��i����e�V{��y$ K�W=�]$�^;�؍MڭIv��gv�Aw����|��)8;�uS�@60A£�JD��xЁ^�̠��v���⣯N�r�L53�p�n���1m�Q�}N�/�J)���`���f*o�$��W*��"�e��Ʒr�/�o	��Î�-$d��]2Q	�M��Wm�� �$��˰��E��g2K�4���p��w�Ɔ{Y�b��q�ƹ�貆bq�8PA���jX��l�`[Y��v�!^�c�r�$,�dZ\��Ҽ�Y���G����+��z�m��Ų�ݏ�`��?!�|�0e���ݬY�R�5oPn��2�-s`ފ�"�B��Y�@%��9��ﴲ@
��J�/D��dj�#Ճ7�N�n�{��|A+h�OзFfU�ρڍ<=O|Y�Y���1���Ծ̝��jd��K��Il�<�W��1!�_L��>n��h�E�^9THo��&b:D��ј�-_F�����|`U[�����SLX�z`�nx�4�z7G^���R�6��#�1=
�˺5D�4}�� ����������ͬ��vK:/8��<v�:��e���K�ԃ/�#�%�@����W�tКq��k�c�/Y����z֎��KA%Nr4�2d��1ʩ���~�y�JK��e�-�z8�|v�x�˻">�%����E0���wu}@G��u����X�B�a/|�E|[�:FG���lr#}��HqL����0��{Xw#+3q���=@�"Ѐ�bӭeH�x���Mo���,��`q#��OB�[��s�O��#h �Ӛl�DE���SJdb����M�:rj�("�#u^���[U���!
݌3��h��炗����`;ص�IӇ�l������j7Fb3�Yd��_���
Ӥ�5\�I�YUٟ[��[�����������J�Ϳ�&� ��L�;=��f���	��m:@��g�!������	��k�.Y��������મ��bi���$�C�CQp�_��l��K��Z{�d��rW���6f��zރk�~fA=͙���z�{�ֽX�/ l��uK=J�j5v���V�vA>)�Gꨨ��6؅��m��ȫ4�?��6�8����[��Ӌ�y	� ]ɰ���)]>�����*��*�6�+	����YT���o@����t(~g�C�0n���@����=��5,��AF�
W�-�ѓ���M�1dm���9���m�{�]��1�+��)�����q@2��V���w���(q9gGӆ�����=�wׂ_��<�*k��z���aQi�M�R��չ�m�78b�3 �L����ɤ�,HX��vWE��;����)#xg̠g�>�~�O��s�H�)�^�J�� 0-{�?QOf>�9s��'���mL�qV\W6�P$,�$<۳�vA#�S�����,��k����v�;¥wWc��y'&6~���;.��ssl �-Ud_A�j܀E]���*3�>o���� ���j^�,.�T���G(�VȎ��:G/rg� ��=o����w���>Yl/]�8ܮ����/��	��K�T��T�/�߱���`��&�vC-�{�G�'�'y�P�fSU�/�`:˖�/h<��v�۴��X\���'%�A�!��� l���b�j݆l6�>g����A���8%�sw'�8ip��&;�'�[��6����A�[�G�| 
F0�tY�je��,N޸�B��rI*j=�{�f�2�jV<�r�O�Ԅ�?�f=)�A�V��?�4�B�5Y|2�>�Jgy�㐈��'΀[�<U��N;������|�������7����ޮb�jCGMU� ����Үd�6!�(G�Oq����מ��>C��<�$�ǹ��Y~�)j�%85��eE�L�L���a[�3So����Z�����]+E�k��aJ�������6#�y���ؚ�~g{[B++��R�˅S����{���h�g�ѱ�%ۥ�لF�h��?���X�[�����bp���}�!�3�?}2�W��@9�m��}i,A��,�j�>��,�]bc~I]}�j�>��p�[�G�jD,o-�o�PmAŢ��(�mP�;؜V�ߴ'�m��G�j��j�GȺۚ*�i��Ե��L�!#6g]�p��Ji����mԡ��J�[�(�A+���[�W`�/��8h�u�R+�5�`oLʴ��pĂ.T��qc6����-�*��׷GeQT�L�/Jw������FynX��e^�{��k���������ɿ�}�v@�;cs&I���E��eo7]���##&!q��'<s3��A ���p�x� F��YSVT�� ����[�J�xθ?3��g�p�6�"S��(���Xy��(���7�l�Yg��������~w� �z�d��α�ۀ�~<��'�}��G�@��!��8
"��.�=�B.�#�R�Zs���d�NZr`�Ma�'��+��=���V�Ӎ��������������d^_�Uc/t���h��(l����DO1�+Q��ȶ^��1D��f��(O�{q�R_J��сw�9�?����~ �»j�8c�&z����23c�	
N���ͼx��w��w����g�hJ����#3K@[O>*�~��\�X��-�y�����X�QOQ.#:n�~�$�A�*��N��8�$!��{�&(ȎF�O��C���R�j!��![,*+3��p�b�l�J�\@L�ܺ鼎}���W4ovN#�����fƓ��x8t�4�y������|n������&��,R?������o|�����)��K�Jv�/�Jr�� �*����=� ��ʶ�|��t&����5geÛ�)8�ozi���U9�e#U���k��	F�:�2�@�?Lv`�6�(�3�d���6�	b]��_�N�^+�~W4����[��d[��k�K���A񛢊\��%�A:anV�F�+$j{*ī�<���|�nq�����xl5$(�q������w{3��'n��V[Kl���c����E���%�*���M�y������s2jmhT�*F�M@}4�s�,`{���gr��u[/�}i_�L��j��-�	����+�=W��y;��fE�_uձ��/��j�&�����w:���,[����pBL�J��7oꞕ�,0��)J�Ur�\���_��LL �a��}��|�~���T��#M��
�{ݸ6�\��$qJ�a%͌�gV�3�7 ����`�D@bhrg�A�ï+X���d5��āiه�hT�R�q���i���8����RS�{N��ϧ��*B�I�r_ayf�>�)�I�D��2���z�ed��/ŲcH���m��O�@Yye���I�|{��C�����y�b�3�\w�'�z�D
܌>S���h���������7>y�����dF�B�z����W��csMoZ�U����Y�O���@0���K8|?=t2�>J��? 2.	�Fa��ך�A�ǜ�{>_���|A_��1b&8�������8��b��&JF���n�ĕ�l�&7��WLRߙ[wɜ̰�ژah��!,zõ@[�4��8���H��~Bz*���}�������Yr	�������yqYyƱ��D��"�pƦ;�8�I~Kkf�f�B��C��3]��vw��CF��u �j�B@0g�n�C�e �J��h��'&�����W��%v���:�Β��S{HwX�Fѡj�:=��AS^�U�4���w��@y���QQ��pL��Ʈw��3��癵����ucGv��bх�@�&����9� WLC�Q��9�Rڬf!j��c |m8&��i���9?���[e�>�Q�V7"޲ٔ,���<쑳@fޅ�(����5Aب�'�����@AvW����O
���E��h࡙��O`
��Ξ�f��R;�'��VH�Z��Ȱ�B;�j�E����7j�g��V� �,�
���#D�b�P���刨psݏ����乿������CʳS:6h��K=yᱜ����6dO�txǵ��� m�Wi���.P��cA�ؖKïK��$!��\�X���2�{��l�~��}
�[�<�%�?���G�9�C
V�9gn+�]���H�bσ��Z�餀�X�Y	�H	v���J\�����J�s0��3��LTݔ4v���<��l��f"�F��t�JO��qi�����SC�:�]���=V|62_�"�#�ƥnSV�y�6�(�7�D/��k�<#!j:L*�?�vw:k���qt���.-Ddk+���E_�l��VQDS$�KH��#;�Pҥ��]��7A9I>C3��R+e�*�Ds�=��bۮ���m�ь-:�i���w!��ND�p[7����T��.8	�#⽋����
bp��T,���$� #�7FC�q{f����ܶx^	I�K��L���6�a���_p��Ba��X�iM�k��Zmp�q!�g�`�LX�Ǵ��9�y�y��������q�?�Bd�n/l���:�KjF_�!�|=x��3�@5"Ӵ����Kg��qp�eUs� /$���C9��a{� 3O�H"���c�p�O����t������Sh���X��ii�cצ̊Ot&%3%m���*^)C#�tE�;���Z���gk���6J���)Yz0�4�T��9�9|G����?��6�P٢��n���{"��V�	��*ΰ�5�&������h�2D'���������8.ER���>��G������YlF�Ͽ�3�V�4G]=c�u��ARR��I����M).�EaȪB9 ����4-wvp�#n���o�Q����z(�H�낏��:����[/ϝ����fF�u�
i��5�}�4i�l�`�z��&gs��	�V���E����Dp��"�l�%uK�g��z`�c��v��Z�
:��b{�*�7]�ݡ	G�5v:�����i�#
�x�-C,�F��=)7�yӦƖ5��{R`�o/�	�d���o8m�_����6ۃ���s��ym$�R����j!�6 {�D,ٶQ�glOA�(�]���P�	(�j��z�s�P反�\��aˣC�E�Y'�:P[ф���xd5�f��k�v��:����`�?���e<2H-�j�����Q�&Xh�oќ5�֘��~_�v�&��	R���r��J$�;�ۑ��ZVx(�X|$J�/�c�����%=����tK��-���r�szCĒ=9W#��HW'SB>ӌZ�#����0��>?��G�!�rFҿ�.��$�v\��&�-��c���� Ē�U�������Sގ�����D7gY��;�
:�dg���巣G���a���4�a�v1�r��c�L$��^��Ga�_�[���[�m��F�3^nۉ��	�g��u#9ݩ���x~9x7sf-�xD��T�*o^�O��B]�Sg�T�>6�W֚%2A�֯Iٛ��l�X�^��V�C�#�Ո�ث�3s9m��Բ����h8O�Ւj���gJ���0�I�\YlEH�j�S��b�D��9P�
�yb-��r�m��B�I��l���;ߑ$�`�*�OM�	�+�h��'��ᎫC�h��-/�N:̑o���tT��'aUx>)\C��f�`��C�^�^����y��T�\���5���B��K�nb5ZV�g+�F!���}�h5�u�0:n񞉖�����$0_L�j�R�ujK\勽�Z��?�Z�/?�vJ&�����M&�g>k�y]��aa�b���l:=z��(
$Y�����73v���n�\YcA36C+���@�\�KC�{��[��^(�S��A wZ2gG�0=G!m\H�I�����=��AaVl�cey��?۔��74����O�l�~֠Z!�C��Ǳ���#�,�K'P��������=�֒�X��9Q���s}"&!��%�0b�m���M�Y(=|��O�äH�\�=嵶+&�������ܟ�-�,6 t��^��E3�*�<�b�����Yb���;2��V�\�b����\ɹ��z_��
�̬�q���f�� 4lZ3: 7n'E�me������]��jI ��/��^�mm`��m�H�8�kW�#hL~c������L��i�I�o>H���^P�j��_{��-0i��{�QGl�-���H��.q���vMq��"�%z$�����I"?��c� J'K�S�.�"!�e�+�t�n�nJ�I����e�Ғʪ�C�w��5�h�*ߦ�2��X��$T!MaI��L���:k]�ζ�%��Rh�I0�mm�qc�f�-��Q舷�ܡڈ魌oV�ܘ �}��d�7����)s<�Z�E�"J`�7
d�=aD�=���2M�hB����<�,�zG΋������.�2�Dm�fo�$��he]Ա��5&��C�^t���!�#����j*.�/��ݹO��T=�N6���]�N���ķH~�`�^;���5]M�j�Yo�e2�(YӚ3���H�����@����pw���/��)�h�L�������2ӣ�r��Ӌ�q�i���e��>���@$�����A�|���[��������=.qD'��l��2��g�Ro�k��/c�����[���49���W����\�CݎYi�m�~i��DCGxJ��N�Vcډ�٤�?���Q�P�e�2����o�S��t�R�H�A��ծ�7���R�a�ޑ�Y���v7
^&�޻r淍�������nŵ��n��T	�B}��+	�rk��+I
��>N݁]M�w�k8f;���ǁBK��g���P;��HGy�-'�a\)��z��݅�d9���J�~4/p�J�Lt-�B8���&N�?�C��1UN����(Bh�n���詤l���:�@6J�oZ _���b�#���*���6IZx�����_򪬪]�9�F�PF�lP �א�W��(���1����)�1Er,�xL��]2��t���=�Ͱ&�Z�O��n��fJ0��|�N8�Kރ�GeI����� =t��! 5[�΂%Ɉ��}m��1]��U0/ ܩ�T�1��*L6XT,��c�~� ���F�9Ĝ��:�t�̀��P@î�!��g`4��}k�# *��6���`��Z֫h����u?��٬���Myﰶu��'q<�_#؂�P7���𱹑24/��it��u�r&�RU�l��A1���؇�ib윹,J��ԎJZwk]yf�S�1O�F�<B�C3��W�à��|g��e�ֿ�+�z�Y_	I�E��}�W���X�,5�&�(��g���m�z��nMr_��]U�O��;<X�
Q��*8�ܰ/��W(�x�����T�fB��82��!��ne��q�3�~�vG
PHx?��'T&"Ҭ�.l�E�Dj��7M���^���=/�=�ʗH������ٚ�6�ʦ�?�� �w��E2.�).��Vu72,5�+�i���;.��z��w&�?�0��/��<�4do�[:�1U1�І�s�v	����Dr,g<U!����A��"S��_���?����^X��N"�F^r�I���.w��@h�����#ɋ�*)|�q/jwD��|sQӁ��
rvmx9��K��	�٬����R��J!�Zmkɷ@to�s�?J��$�f�~�)����<�HRuJ�)'WMp�)\�e܏�����f\��x ��E9!��7�V�����R.�hcwc�tN N�c��!sJk*��{t����?�}�>]����ć4P�ٖ�u5�����h�	O��z7r/��|I5�E�F.���0ѳ�	pyg��y?W��9��>����!H!�"R	�)���7m�� ��Vyȍ
^:�WO�q�[J��z^W��D�#ʷɃ�شʬ�t���2�s�]Ym&k���|K�.�gӆ'#��W����n��r��d�wS�C ����mB���$djVM�h�k��+Kf��w��̉
�3G�9���<;%�(1�0ؽ8M%ӣ�=�\"����3��G_�(��Q>��ʿ�����O�䃎�J�P��(�qkR�^>�X`��Y@N�5��r��.!���9�P��ԾΚ�� Z]��"([Z�CS@��7H���?f������=�{�'Se�|����m�\Q�sQ�6���B�-#��x�l�a^@�V��J�����rf��:̱K@������j��`����w�̎��y��z�'kZ�r�G�����<�Ȍee[f3<�d?��N��B��'��@�ʖ}g���|M]\x�V�Nz��s�kR�Y��`Wh)ED���QN�6�К`�YS�
�i�&�К�T��Cx� ��آ$6-��*:�à��73�����ٔ��w���m�g&�QPdO��(�ˤ�Rg�����Ya�`6x�K�1Eu,�,0���^Ll�%��)���#z�<?+�t��0)^N�y=�|A�ՅM�#Do�)�Y������r��WO��D�]>�d}��o;��cQE&��}Ǔ-)zi��<8�w���M�@G~�[�?��?�$�0H�-�\Y��C�pϠ #�t�a����Ǽ���wn�i~R9 �rj�W�n�+Y�>3>;��-2C�y��Z��T�<��<�ގz�X��J���H�`��\c���I��T��m�?~taLŞ5��ɡ������k�M�A���4$��݁g�
կ�*&�
�0��]��������{�[2��ϝlXh�N�zES��6�msR]�T3��ŝ�	t�@���e�����u�RW��� �I���,�R�j�C�;��P��a.dQ9" ������{z[ZXX��p�'̖b~���_CW+_�������FX�������ͳ*M��:s��Cq�jh��*>S�z=*'Υ�&+OG%��{��N���[�4�L�-�?O�|�Oh�Ơ��a�-YҬ�Ү����>�>"��s��1��ĕ%�txAf�i/;��T�KP X��.cl[>K��衡1�+�<-8g�5e�=��[&H�����u¿�~ ���/�_�m���)���$];���އ��c�s�i�C�w�^J�|���[�Z�٦���Ⱥ�	Z!։�e���1�#��Bep8Z�I�t}O��qw�hK�,�(�{� ���\����Pq�s7����-W��GE��LI��^�IP�K<�w5�x�Џ��Ιz"���+-=���� �|4L��3WP,gq�GW��	_b���R3��?.O�]a9_t�M}H���H���ш̹$�N��&��������K�9�ӗ(	�}��	�-�C_�Ja�z�r,�v{�B���w�%2��w�)�vf��u˕�Dx#�(k�L:4��{y�g�s|t�w�=��=V|F�c��0z���,�>�35n͔.g��g�Q�Xq��4�X}�������k;��/�{�V������i�jWtu0��7� x�,h�6���E����������TEG^���7�Z�����F�����t��M��&��0�@��P��k{�[��lf[�̞n��z��m=@��e��
a:ݪ���F�D��j�&Z�����\˲[Ai�V�Ǥ���
�	��mE��\k���ݠ=���:y� r�د�L�XX���Um����|CC�q�XH���o�����({���9-�B�lJ�"bJ9"�:)f˔��#L(/���Oz�F�d������!I� �*�Y�@ ���O�<�B���A.)�bP�(�x��:�"��M�8�2���Hk�27��?dw�$�TI���c<sN	��w�����M���$��dׅ|��p��;��:rwN���N�9[�!��A��{��<�hSD��W3
s�x*G��	v����1����tƩ��|!~ӐN���1b�ʑ��m��%��Rs��}y�ү�Ůȋ��r�#(����<L��5�Ǉˈ���)[��J��hP�[��]�2o��֥"�~Ě�Tl)���h!�ث�L2A^�.�(�b�����H�+g���zE,'"( ��[F�@J#a�q�lRd�'/¯Mܟ���wy�GB�X����1�ѧeTl]͞�j@Ľ9/�,#��A���n��>rލ���:�R�e8p:P��N�[e���"�����������L暘0�o�P�pպ��U�=�Fa`A*�o*����4�O��I�|F&ܸ:��W(���SUIz��n�QFԀ~u��6�b��I�7�0���(�ҁ�ST�}�M�܍J�RB�zcܣWJc��s!���.&`��@s=��]�W�E�(�����)Xg��<�鎃r;	�b���}�byRY�XF��!��b7|)�w�E�]%6+�}���
�=�;�L
�bL[v��<�ށh�ӫSP���ٚ2��[/���Cw�/p�^%�E��9��89"�m\�R�eBE���D
���,9����B!we�T^�p8?�.��*R�]g4��m����2��3Z�H��w��<��H��	�wx��v���{VI�9���"΅f���W����؛n�$�y׎g]o~� 
d3��&�{�����GS__v/���ZJ��U�5�*�Үϛ���`H���:=�kzj�Ji[*�3���Jj�cX~h�,q�:τj�B�-?֠H��v�A��o"/T��c��d�+U4B��lPwrw3㇕�6�섏�1�@>�����8J���;�Q�Ur^��n��&ɖ 7�uP� S�f�$MHnfj �&��΍�&H�rQM�����G'�r��^k�'V���r�q�Ү���*�_���;%�^⿊S�\ǋ*D�|�3�3�����.b3~bx$}4�b|;1�\�^��������.�}k�Ű��6* �F�*e����r�p�I�q�á#D3maV
د<��p@ [�]�,֮|�
�]��]=��%���D�{��Ȟx%䩄v�zE[��Y�è	�x�_zސ?��EK��"�ˬ��}ѧTU���D-;.=���	듥u��ja�`z��z]q�#T�&�M��j���*v���<I*�O��%�k����"��Ѝ�Õ�:Φ^;�!���T���v�K�m�%���}��)n