��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&q$�7s-u���Rf�2�F���yS��`s[Js�&/�rR���C���C#���h���w����\L��M
�aҏ�ň�E���h��ÿ3��[�c3{�B�ʎl���.Ӣ���G��e�D�h ������p��O$s�Q�щF���̙����5V2:��W	�`��n깃�"[��ΕvlB���
4X����q"z�7'�����Mxm�J4o�A�*)���5���/��œ��].F��Z�̚����,3�]R "T* �a�B���(g��Ņ�Rݐgyp�v¶6�� �J����G�/T�D�=�`Ϫ��z[�� �<�]��Z��W��r #��]��rz�ag*p}o�q�r����ՙ��H�'HՀ��d}m��<�sf��u��v�H���Z�;�{ 7?�mũ�H���(�=<����r�D+:����f��g�,x";'���gf���B �����1�� Jˊ	E�,��?�_�C7׸�f��Ӊ�A-���,,�U�Ik����}T~d46�OQ��i
��S�g���N?ø/��JG&�!�Nߔ���T�P�"�,"��n�Ȩ�^܄�����&F`{��R��έ���y��D^�Q+ZJ[9<��T2��娋(�+���O�.���	2c�ŋ²o��55py�`�B���VYG��%e9 I���v��ڞI�pJ��ka�y��p@ �8�C��A�?�Ӹ����ԩ�Ǖv1r��Z]!��9��A)IX'>��e�|?�8,uR��bh�2o(\��R��kj%H@�y!5��G����`��rS��Ny�-�p��S�M����ې��@����~�4���@�ךV�D�Z����#������o�8+v�`:��Ϝ��/�S
��cFM�e�l�,��[�޲~��Ă�����K�p��E�e�*�9�mɻ�_hEW���d=	��(}���[�k��l`�n�S��$Ɏhh��徸���$��t���O!�@�,9�E��m����ET�_��D)�ʐҜlU�9l�F���Ȕ�Ep�4��þ'�-=��ؾ�X��-.��ns!,�F�'��FD���W�����e��F�7?iΉ�ӎ�^Ez�еUF{.��HEBy��Q�젹�42#��/gF��kYu�M5�q,��ӎM}����z���3�n�9�^G���T�-X'(c���]��"�խ"X�>;\��YE�^����zE1�u����m����}������Zg;��Er|m�Y	�`a�80����y�Մ,M�$:�|���>*�ƲTA�c]75O�����x�f�Z\�Z$���T�l�6Ҁ�CO�i)�W�.%���@cg�|S[�N��H��d����L��'�G܈���>�����-mElE��1P��re�f"���
�:��S�J!ƞ�1�N�:�� ���O>�d֭����:��EZ��lW��
Nz��޳�܀cT���yJ)�����e�����Lx��o+����6�)�:�L,���|�!wC�9QI�*��R�3��,�uM�����P�KZ)=6����(\�[���Nf�Q�\z��݉�����ǽ�EoF�"��۱��x�&��5Z�}n(�!�1�K��h�h�<��+��Ōic3�Y 0������,�-[)
Ԟ�=R�1
#���<�~�087&��o��.�x�d��;�{�(DI���D�5s(�Hx���_�C��ͻ;��F#�2M��hk-�Q�>�6(PM���K^!)�c�HJ�c.�ʵY�2<� �#߽B��n�U��R�g��r��RaQl$ֆ"�Tz��Jp�Ԋn<��U?�h�Q$�c�O��J���cjK�G��@�J���Ĺ�:k��;��[3��w�tʁ�,U���M�������ɱ�8����^x3e��_j�≆���N�����q`.d��������c�Y���e)���|����}U��P���uK���ֳh��̃^鞍8 6�U/���(��0�����{�vU���ت�r<�>�2�oU�ӕ��\��3I�X*ů\]P;�1u�}e�Jq��w�<��-��K{O����=]�C^�J��U^��b9|@��b֎cI���s��ʕ��&q��G$�0ݖ� �uL��^������z�qK�O��2�t��MˎĻ� �t��������)8�._���ؔږ�SL|�b�bݰSC�h���<��wK�z���sjXoK �+r�W�G
���c&�*@��%�C��]<z\����a�����^��f���U��$����ɸyNDG/�'����^Q2s�r"��=�RKA8�W��r"	�3���JBX�&m�ևt���uˁ �+�d 1�*���]��N����8�π5Y������=��g�(�Q�!�)��"���p3��#(��udLi|Y��LŞ�+xG�� �S%q"#���LT�p9�������F�����P�>�rG�_�(	UxKښ>�kI��e�)����xl���[!+
;�^*�:�z7���_�9�S���e����1=��\�{��0� �fF�g ���W�ߣ�Jc_{w��(���(]y5� ,����g`R$��ե�ղ�G���)����pn���s��������\�@)R�}�,�L��7]�{̈X��QC����)�cIF��5rY��)�7�~(�6V�:�ĕ���(�8P�嬏�͖�#�X�5;d0���@Q��,�M�P7�qQ�b�3d<�G2��X������|�4E�xn,�a����u���DAe8��U�B8�S��� )�^�O�	.��G�U��D����^+��7FSp����X����Ȣ�h�����'���+��� ���L��T��0�A�F�/e1�����p�8,T Q����g ����E;
�G���k���0�cb� z�;�9��Ê�]���$�����6;���iW�ՈF���;#��Av���NP ���8Y����E��'ˠ�Z_a�{�<~�2�{��ߡ����T57�X�[Y�J�NH����9���!Mބ�Xj���@��%�ӻ\#�a���@�_D;�u�b�AL~t5�;/�4\���4
�MbٕmH)����Sz����3�nP4_��b�K���󯻜e��~���ݯh��9|��>e=���L��u��_�+J�^@tԁ7W�C6�W�|8��(rT�٨�A���hUUe��X7zA��{[�	�)�SC]���>J��X�1�4@��cw'8X�t�/:�9/�B+��`���Ł0 g����=5�g�pl.&��$Y_�Y�/��j�����v1�5-�������Ռ����ծh�T���4���eR��̫&װ��\���Ң��"t��#�BH�D5�
a�Q������Y]Ն�Xi�~Վ�2�=�'I5��7M�;\��v�
�V9�涑wB�iгJ�s�`��)����'ި�L�buǂlxE��lz*^B���%���6���q��j9�+Ķ){�^�Rqu����	y���@bV1V}�*�s�xR�ȫ�J7V�����O|��l���}���ڰ��Ro �ͱq&t�`�|@g3�n��G��i\Q��r�č �'�p"e	���ŕ�����{�N?��0P��n�	f{ʨ��U
F����A���JݖpX��k'�1���@)��l��3�'i��]"��>���F@���q���-U/���NDEo��߀��y������9Ɠ^�tQCRB�{ue)C������i�/q�*⏲�/����Q�Kc� ��_��s�� 6�2�����戱�W�Ȗ��aƔL_̨�B���I������ʂݱW���!2�$��B�����UMM�����%�7�h[À|��es҇ǁ\��/�Rw�*�z�L�YMڏvhK^\d`����ɮ	|�.�ͻ��Q�Z%Uzl�k�[Lbx�o ��(�;����'�*�)���j�B��<�-�匞T!e�R|��=!�8@��p����S�P����^�	�i�+�`�����P�iO��%�04��l���B]�����|��� *�px��W��`�"���������*4����r�-�]o��4B�~��3E H'S�|�R,ȇ8c����ˆ�/2�,� ����:,u��5��qlDK9AمPi�b��yBk��p>����wo�txh����*m��N�<Eh�ᗲp?X����ʁ�m��xN�q�l�0�� �N�a�3L���f�˸T�)��B`
��pt2܇8]僞�JA|]x:�p1�;]b"Ej���� t�BxC!�Z�'���i����(;��_��q�s��B����`����RxX
���q�����Is�x��쪼�at@�.c���:�܁�SS2��s)M�Y�+�]��h�E�a Z��8 �s��a�A6��yx�TZe����Ѵ�Ƃ�GP��I�B8�a*a�m:�D��'�~$V=c����	��̅e��lA!��`ow�MB$�+���4¢J��[��Z�t����@k�]3\oǔTY\�x�4�}_�Y��`l�h� 5��z�#� d�݋\���8�k�T@u;�3���/��>�e!����Q�ǄҘ���B4&�9Ӥ̲��[>���O�q��n�������u�m���D4�Ҳ  ��v�m0�YB!Yz��lP�6������[����#N|��p`�i��*
��/�6pM��"�+�K�}�N�w겫��q�B��ܒY���PD6�i��y�o>�\D�>�!�T)/�C���!�V��X��?i�3]�jpf��xy���|Ć~��u�(���;��/��2�W�h�!ze�j-5lD��=J*K!�؆T$IHσ*@�� �IQL��q�!q��5��d��1x�g�Y�~��Cg����3��E���)�^����˫˵�FL �d��3��H��M��U��W�\�{����@_�/��^ХZ�1o�����&hz�}����+���F��x��� QA�#� �C��v��D�=�͹5t�(�� �G�q��0J}1�(��ʧn�t(OC�*Ř[������c/�% ȵQN���Q��|&9�u]o���	u���/�7�#��ddp{�ǘ�:S�y�(OAG4�B��S��5��"'t?@�+�ef��A��kX-���W��Ll�Y�"��ܔ�IJ@ <�MYl��pts��n��G�b���ee�"j;Q�%㖟�oA&J��-S�ij�6Ҹg�'��8B�&Oa�Z:L�Q�����M�=��x��g�+����e�hQ8�}~�ݼI�G��!fA6ܣ��z�zw���ϐb'�Z�������߼+���)������\H"���c6`-����`~x��y�ZO� ~p��M:0SçS�|��EE�߻}�$�O[P���T��sp.?�xğ!�������;��xz�(m��q��q�-�u�c�Zը\�1����e�UE缝6S��^�f�?�"{H�{M�ep�B=�\�U��n���T:f�~����˘i��OGǼQȑ����Y� �V74��#�(�W:,��f�e6�*��_
�v�.�"U^�' Dl�#�xZ��)����c� �s���[����'QU�VH�6�K�/x�+ؒ<�������Rs2rv��{�?����w�Ħ�q�?��,�GT\�Lی釙��_�A����G����Lk�,-Zl��ϕ��PdĿ��B5w�$��m�]h���~��B���b,�� ��#U�x��^�Ju��m8f��u�>�S 0	/pV��%0�����Ƴ�o�;� �$hC�n�Tn���hS]�Ԯ{y��,�ICQ>T�Q�~�d�b}�u�Xk�;���Fo�7���z�{MWW�{���Y�d8A��T�ֻ�IRGwI�:¤$6��.��s8����\�@U�en�g�U:���y���:�Us�6f(LSç�#q�m�!�d]��qQ��[ ��$'@�'�C�dv�|�3���`�{���j�}*h	O�%��#����TP�:*�&�����3���f�d�:`��Z]����I�~f���NJ����D�O0�{��iw���b���矽ʲ���t,�~��,��ު�qѪg����T9}�ƿ7�Ɗ���Bo�N�[^~�I>�-��W�> ��s{- ���(0
b ���LF�p���l�k�u���n!�E��xP1�eԴ�y234�M�\���|U�Fq7w�6+�`���d�{��h���(��T�k�B㶻�4b1�*�����]L9�����ϰ��AS��uV*�y�&e>�!m��ՂO��_�L���l��ӈV���!, �B;�F��?7o��]�k����ؽ��(d�w~�>��~�n�����+¹�L� �׸�Ǵy����f���z���7�҉�����~o"n<��?��g���n�?�����k>�b����2�' ��"	C����]��x]��(F�`w���U	x�x��wD�d�A���ib�[��E��-���q�L��HJ����\ۦ���_��C,>�p;��iJ���żàKӘ"C�� �Ԕ� �KA/���d����M����a��J�.�ؿ�orpMp3,i��y��H��Gh�W��L�i�M����6�#�Xa�c�yƥ���Ĳ(��u�p��ѽ[��Rs8>�v.P��y�R�F����`�}�G�F^*�N_\bʞJͩ��f���䩪5OG�#�>k���V�e@�]��e:� �{��
��Z�\:;�xd���pa?6���W�_�R� �� �8C���^ߋ�?G{|+�A!����/ŷrke�u:��@rj@����E�؏��%����E���~�5���h�S�h�ɠ���5�D��儧��cV�k,n�P8�W5
�	X�>���J*Ω�g�8l�aj-�ۍ�閭@95U���^�8�P�*Is�<�;%��* i&ʧ�HY�¼�P��Z%/*5oi=�	�2��)D�E�C����_��m��,�3{�Ry*��?���&p��V.�,��9u��Xd\���D7��Иq�4z:���m����z��:�9iW��)%)2t�Ơ@�Ϗ�$��/����Ή���Bv�	3��>C�$L�/Q3'���|cbH������]��� ��Mm�����,2���4���mv�����c^�#�����%�:��*$0�)� !�� #�!��pw�*���_�M�t�~��#�4�W8#����W�����n��ƗH+���g(W�A��q��m]d=N��bQ[�M�=r�~��.�b��y�N�v(�Y �q�nP��(/]�9��.��[׬�鋽�^���$�+�!W���Un��R�e16éؤ��<$���Ed0�t��������$���9�A!�,�Up������V=� �,'��.�2���=�W�ɥ}$��hh�?�.��o�j���!f�qM�j5]�Q�H�������
n`xôE'@�{�-د�W!�Ud�_VI�q�����8|�Api//�Lq_�	`�oؼ�>�.�;Q$�*S��=�հ̞����yW�̀.;��u�]�K���{>�ݦ�+ t�S��U���@��aA�������#�H"���-=g͢��ʎ)tA��G��������Ji�9ALS�2ل��Z�w��
�s�eoI(��;b�o���&����UJ�!	29(��^j0�q�n2hS'��U�v���A�F�٦1�'ލ�Z�iJ�	yP;!�A�0ǟb��&��j��(��5\i�U�9u>
J�>zU������wg����.L�o�9�:�}:��eP�O�H5:�T�bV��Ǉ��-�-ϭ ��t��d�H��9��%��1'���:O��i�c�K6�m�-��A�i�Df)D��5ʦ����B��8�� ׼v���ւL�`U�l=�N5�)��__���N܊���+X��N�����&�$�2�����*WG���ͳ�f����2���t�gg��a*�#P�q�[q�(h1 LZ��\��pW*"ۚ���զو�GI�X��
2+n���=
؞�=�.8Q7�3�#������Y���a+�������?�eᾱ��I�#���G�k���<��eQRm�*a��v�����>���T����6:wi����3RZ?MW}�T��� �8@)�_� נ�L�����sL�a�0�k�#}��#�����vg�%�[NLFu�'�Hq	f� ݰ����),�ǻW��a]��l�DgC*V�\����Dwq�Y��_Jc�rϱ����7�T�F�XmrȌ�~�ùǃ�x�%懄��8�i����\e����� t��.7^v�i��	DZ{z�	Coo�������@���
�0#�v췾2��]���:��)��[J�s�|����iB`���;3��7����N@�)C��eD�ÈUM	@q�,�yBi��I~1kV�Pegȵ�	ԝ�����_q?^H��Wq5-�_YU�Q�EfP��
K�Ds�X�[��M���/�*v�g�zu?3o�`Ϯ�P=Ŗ��^��E��2�?}��H��<���~E�0�Ϸ@�:+�hg�,W` ��`�MIQ��b�~p�%N�I	w���*���t��=mL=�ǮUXp�j,�/psc
&�$�9�LE@�4ַ�7�K:��f7 C�0~����]��Ɇ�j�� A."&_����$��?"��/[�W>�9�گ���p��>,˝����Eݩo�T���ݥlE02J1�#}�Ł�^��M˜�6������y~r"�5h�\���i(F�8��De�X�i�Si��A@�g�}�i��>e�Zq�8{5�O��"�0�7C}N�z��Pe�T�E������ئ���9B��cKoI��b���/�u�dZ�#o���$�I[wV2n�0p����I �>o��/]�=.�"����ҍz<0D	��6*"L?<E
���S�2AM�'r iV��e7�sD�r6w�b�lOqq�*�1� z�!E{�p� �<�V�{��锁�"B:�~�����c.9t�Q:�	x��[r��g&dt���/���X �KfBx�M��H:쀰mu�ډ�o,%�d~2�(&($R }T�t��k=tC�(�_�	����3��S��q�V�Xˁ����w� ��Y�lT�%�"�G����_H*n��0v����^�R�9��j����.r\��B4�E���&�fޔց#,�!ED�T�J�j��#�uSF2�HcM��Y͠9f�o5g2/���um���ER��`u��b���J9�[p]$���{˅�{�� P������+�Ǿ_'����:cv�������N�jF@�ގ���C(Mۿ���}��`� Sd���dT3!D�̔>���-G���մ{�8;2V���-���gs;�6C"}J�[�g��� �Z����e�u|�~��2�̐�E-[�Vw�O,۰�ڮ=�Q=����$��!��#X��ASt�}$��zm�R��>\)=i,I@K�n��.q�ė����M��L$T�.�����cҭ�aI���Wr �� �7ǣ�i��-ƅ��Q�=��:��A4��.fPkN��H]�W���/K9�1�K!���,�Zh���a�>%��᢮�5?R��6Fiup���x)>L|���!C���me�/����;\�#���
�DD��S*LO��&~[<eqr�I������h:?#��I��(��Om���?�o1ZW��|68wXH���׳��+�ʫP�i�#���1z,冞
�"@8��E#�?}����BR//}��ԫ��V���=aru<���M��dH0ݙ�mdұ1��M|R��Jۀ�U(�5/��l�'0�Vj���ˢ��Sӕ�%"��#�7�Gz��hi�վ�Ҁ�xH�ʂc����T|V���X����?���zP�@_��vX�D���]W?Z��Q�vvd-�,�;S�8�UQ��.�4NH���B#E�8��(cHͯM%(� a��,���$��p���g�5��TY5����aNd�L�|��Ζc��(�)��1է�N�?�LG�È.^���榢��N-���&��a'�ޕ䳀�Zi����p�����w�� ��&�_<515:gZ�ا�Kª�6�_� A9�?ֻ�"�)����.L���|A���mBm|ݯir��J4֚7K�a�s$?�a>`z�Y�C7����.�Z���N�d؏� ��0[�|g�8�V#�R��im�r�T�Jm��S����Dē|o�ޙ�]5K���-�[m�]7��t�4p.^�,�B6�Cu<I�"w��١䖻�B&���́7�Ĩ�]��~�͓�����O²4O�|
����D(�"�����`�$)��Q�B$�u7���}Cgq��G)���~WZ�B(l�9�(��f+��ޱ�TL�wb�~�����X#
'�p�����A���[+=�����BmH���c+v�W��#ֿ��C�ZO�z
���a���DEZ���0�"�����`S�����qJ�a?�p���o��-����_�~������C�M��//TH�qx�O�0pg��!����J:��^�/�+�����:�p���yCC��C�<��P�,8�_!�VX�����{�(_ٺ ���e���\�f
��Ҕ�~U���)��g���8;<C<]�ž��&�ꆙ���Zm=��⁮ <�G{�4�C]����U%��%��F@5��N�캴���6H9L�1�H�A"P����w�;�|u�'7���7=�i�/�e���AJ�5_�p�@K�������\}�C$l� ���Z%��m:N�i�P��N#m�vn�rn� �nj�[r���T�\,�M� �{�`�#�e���`���bxK����C$Q��d���ފ/`}�Y߯�B����	z�5������m����O=^����uR�4$}�J9��}[��	{�J��]x��k����s��,��i��U���R�����:# �	��v^���$	��){�������6re� k���wA s<�4��XP��x�ݠ�ЃK���-�1�lw�6[��_�M��Q�D}�`�-_�?��u�W]�j��4D}�������ty�g~n�[�RB��]	���[��=t�8R��싇b�{��n1"������y��+�ŷ��if�'0�z)Gh8z�>��!Sx�= �W�\�� 0E�C[�9k�U@"{@��9Z&/�$�\ta����qff�|D�fWsF����*���}��L���0�yDזz���h�^�ݥ�
E��;$��oA�ŗtmԸ��G���#I����f�в���z���o-�++�l�q�̀�)Bt��w bT��-�7��$��w"����� ���i���IJ��88����
em��RX��y.UE�T��cMa�"3ڍ� p|�
�;<�ϣ�.�b�c��U�[��p;�������i���Q��O�-i���`��r�F�D�H5�x������q�����-t�M憓�E�B�r%�o�fKZ��Z�A�:����CyN<�]���a�w��RvU����ɮ��K�n`�d����\.�d#����kn'é�D�
� l�;.
s����2+/:�'	�(T��\"C��o^(�v��"y��ȍ���§��G�[���Gv��(����k 0���Q�F��2����g�ܯ5���2�r=3�:v���^���� ��?��}��Ε҂��Ӑ��ۂ�{6뭒	�%��J/Ts���救:H�a>o!;���ְ��o�Ml\$�.{+$݈��d�����BΓ�D_�lF�?C�G���L�P�c1RXݨ�6_߾���4X�6�`�\ ����j�$�W�v�Q)d��l������K�YZQ�8�-�1O��Eg	�(�,���{��+6��y���5{ƫ+{y���d�v�Ȳ���4�8���x�̍��lׁ��>
Y����_��06�#L�J����� ��>w�����I����3����=�Q�Z����y�#��yQ��
kmZ/����3a;��PD��(��Pj��N��S��s���-���A�����+�ͨ�M�<'O��#a�/�,S[���D�������i�����eϣ��tJ��o552�j��~*E���[Sk�8����2��Ͻ���0�.	^z�+��˫���y��!��H+a�V0s{r�>���k4�wS�l�"k�X�:ɠ��~ɓ�/O}�ꌓ�Cc ��&�7J�A��Q����*#e�y:Χ.ϙ�S����	�Č�4�4�"@�78�c&��{�
�3b�U�
�Y}��J�X�Y�t�O;������Z�ɟ�<��
�Z����b��~��b��֒�'Z������D�6eŐU�gW�ہ��7��R~�d�n�#�,�ݧ 3���@�Mz�K��=�TE�3�(�bA�H
�����^�x"�V�Ip�8B�6��,��D`U�,��5�2a�0��`�C);UL�&��U0�>X�^�छI��	��Q���02�yn�-ŀ�V�g�	�2}� B,R���P}Kh�G�\A;8RZ!%�<"�t�N-����O��Z�c����!�b�%XS�o[8w!F �0�}U�k&��#_emV:o{��si���R���P���_ �����0nyl�
S�)I�?�M����5�
U��"����`?�!���^W��F��� ��F���2�`]�B$����Q���ݝ�6 �Η]6x�8��8�C���C+��<;�?R�(Ӯ@�@���$���1�H	�x�^��Kۦ\2�SJ�l�?����"	+Rl���h��g��I?�. ��$��ع�qE�-��HL� x��k`�Q�t��|d�k+i!&F���e��z�@�e� R=џ���=�&-W\��Ғo���#��82�ϼ;C�
�r^?��H���.X����4k1!5I�d�q�
'�{�7��(�E���V����`I��}�N��E�����#�F���F�i>'��V���],��@V�q£�<�e@��_A�[��� ���M����MK���(N#�o	�.#9>5:��l0�|L1���|i���B��5��N���(��L���-�����̎Z�{b�ƙ:<)�:����"ߦrh>�e���k���Z-K��j�7�ɺ4X�t�=aZ�>G~PڼH�&^�+]�[��uK�r,��ԑ�w1U�#�o~A/�OW L�{�W�Z�/&�F�i�yy�'C���H0B�Y�W�-�! �\AK��[GE	_f�~�[0���dK['%�*&�GFnU�R����i�6b�/����J1kc��-a��0\�S[%
��*����=m�.ZYB�%=ύ+ő[<R�Y@���b*� ɷ�Q ��˩i��W;��_�
��p�A=��J�N����>�Lx�0�G�p������wQ����@E��j!���?������y�ɞ�iQ��CK6U�������-�+�H�̜�l옮��Oы%*뗅tU�CѾ��88������j�}	5��`�%�=i�Vk"����}��x-(��+4�oK��;t�g�:P��Sf6����H�k#?���	A�<U��ِwU���q:+UfZ
�Č	�7�C���^�����t���tne�F6�z�+f΂?��ʩ�������B۲�x���+.��3.C$�RyC�S�[�혟������$8y�!�:�?�L���a`d.h|-��x�Aŗ�� b���z��X
,�:����Vp�� ��>�6�ܓ[x���H5`T��O�\h<vY_���
���w�g���
���ҴA��5d_xr�ᮦ���u��hF�*��W�
-9��JM��R�cB]�s����9:=U	j \�6
aP���(-71d3¤�RuB�I��8h�\�u�\�͎�Џ�oP}����MG�8Bj.��
9�:5G�����qF8�\��U�y�h�f��m�41g�ϭ'W�w(g�*�sB{���D�Y��w�>�)t���ܢQ����4���_�A&�du���u��P)�7�0�ԎP����c�E�A�&Ć D#��]�5��ݑ�i@.ȁ��S���t�̆c%��nO���99cr�z��*%��'3s�m۟�~;@a|�
^�t���y�Dj���1'͆����ч]Erޛ8�j���>{����*��ڕ�i
�2�%��څnQR�
(B�������O�U��KN���L�TeF�H�������{�d�t��MU�į�<yn(�X�X/ز�A�#�W�7��ܠ�>�^�Jb��/f!$��Q[ΧAA�K�ө� ߚ��;�� ,�d�f~���7ks�h#�℧��^�/LGí���S@KE����W,��[�����u��k�#�S������7�: �`����-=���H�����ȸ|DE�(2,Ĳ`B	��Ѹ�"6����=��D����4;��U�f�e�����.�x�6{ʲ�q��f�	�O��]b,��}�x�.))_��x�� ��X�0� z��b���a��
�1 H�Y����y��'� Ѳx��)�| �Bu|�t.�r�]Gǆ��|`e�3Xvr�HX�)��^MB��Ai�RTl��Fo6�E���lm�l���.P!N@� ��[��ͳa���:��f2g���5,7HM����b>hrOډ�Lb�x�s�7���GO�J
����f��	ļ����ѣ�%�	 3�,*M������~���F�vJ�Piq�>�L�foB�[Ǫ�s����U��ɫ�YgR (�X��W�����5�~�+� ����}(���w�`�n��U5ֶ�;��TE2�Uɝ��7�{'4�T�G�d�/��Z�C���_B�0�?�>-V��: ��F�ΐ�G!��{�A1�����֟�У�1��["SĶĻ�ԝ�F=Y�r|w��A~O)lZ4�����H�c�T�^�f��u��)v&�� ��"'sn��s)DD�O,R�1�Ǒ��2��_عg\f���ݷ�G!��^���*/�|��h�e�������v,��:�oj˳��qA�s0妐��?�Pһ��',G�J��^�� 4mL��f���Z{l��yz)�7�2�ۯ�b0�+;"��r�@ُ&���������Lr�:M��a���-��K��:�3����G?AKp6�7xJ�S��pǌ�l��EL���Gk�䃊�1�	�{"8L� x��o��}�P�#�_,���Ϙ ���6ğ�5�E����#�dQM��ݮ_p�}�Hu���y�	���H�d��'�f�C����8���m����LU�B���6%?��W�ә�E_���	[�\���H�qM���ָƜ���"6y���㋡ �%��}6ȅơ;O�AC.�'�����P�^@8uSL�n��FG�\3+an�}�-d$�N�ov�l~����ą�D,�^b��~��D���6�KǛ�&����do0X�iE'��g�Sp����+)�������$C�[�@�w��4l>�˴T���g᠇�=}+������0-]L/��I�����u0���rozjoC����l�L�k"bI�G2��Md����qV0�mё�F)d��֮���2�AWI� �R⋄�ZN��`�,>�{�&������ٳ�:a��Y13e����@��Ӧ&o���^�3�x��NO9a�F��@/��8l���i6hB�J�p9�V��ɲ��� i/u�+��jo��Q��Ɏ��������ZȂCs������T�l'V� ��Q`�mG-��S�f:�O��]�D�9b�$S��a1D)�Ņ��HH�"J��)�3Y��rA��J;}X;r����&g�:��C���#G����\S!6�)�O5`�Ԋ����!���X1���B�?��,�����w�o�(�i����x�qտ۸@���?���G>v��v#w�W��?�����	�ب�����j���Em�8bP0G����a�v��!�Zң��	`H4ݶ�o��5���=���ۛ��qH�3]*�ۈ޹���Πw(���lך�Q$.J��p�y|e�����$L�����B�ԖW�SB��V,^�,�z�_�7��͉ԕw��l�{�E'޳���ݎ�,iF�+�<$V�<��Q1�@�+�wٽlL��խ�%��G�(2U�F@����s��<�j ��@��m��<�~��g��Z0�һ����"�hN���7�g�f����E���Z�I4B�6�5G����~No�(ś3������v���b���`�Z�A����	�I{�s��V~gIH$L���q �n��-���1�{���GX�H䚎T�'ɟW�U��:K�|?��i����_�y�%2Q�g3�^�ķ��~�ۧ�- �ew`L����"�HZ\x,)2�ee�[a�b�3 K.$,�jȨh��)�/)dK��+�0�3l�j��� �4<��_����7KM�`m?i�,Wؘeo>* ��z_~�q�&�i7NAG��H��P��b4�U�Q(젚¾7�ΤO_�������%�!��	3�1��2���������#a�����UeE��c1~��O0El��`�GHɕ�ZdN+έ��!�0m3�S�{���Mm,_��3���q2�9Af�J�3�|U𧸻X�$���̩�f
��� �u��,�� ��K�(`d��Ȇ����ҕ�	ʧtX=�U���÷������̖��V�(r���q�T����8�q6t����&���Ӓ
��^��q�@����L*�^�3v��'����8���$R�r�F��wJ�%�"�j�����J�s�+,�s�>x�����Sn�BiGё2����މ�����pAĭӶ��|�Ryf�'�'|Jj�N(g����f����<���0�v�X3=��t�3K3c��VL��^�h�t�T&��ܙ�cg�rWV��Ŏ���/�ו@��r�f�bq��ڟr�����!�3V�V�~j�U���$V�x���V�P�.'(|z�^�f
�<�$��÷�{9�׫yzF�XӝY�KhB��hW�`�B��L{r��_��/��Ɖ4����	��䑹����ް����
T͝$�`�kFb^�R[U"pXTo�!�Ts��1K���F3�	�U �WV.���&@� ���}��E�M�r�S���-bk��K���#3�t�'}���Ƃ���5?��4E}~����֋������I{����S�O��� 0�vT��RJ7�>J�a$H�Tl��L?�%��r�h��~%���H�L���[v�G6�҉�k��q�gx ��"믚�h�nȾ�^-���8aԀ!t����$Fr�r���W.Q��:(�� ����;�m=i�K���EB|��e�}$��4�������0�G��ͺ�����o^uht�G����%�Q�'LHq<i:T�>�d�1Qy�m�~׌��fE%P��)(�C.y�pBi20�V��g;�I��Ь�.N�T�"�a�4�Oc�/���H�n��3pa�X�/�ө�FIQ�n�����H��4f����}?"[�`~�7�Z�9�����+�b"����.�4�t�m����R6�ھ,�ӂ[�mt��e���Č���-�$���|�BcW�<` �����
Sv�-��75�}�=ic�em��6߽E~j_���A/��J�k���0k藾΋O���K��aP��*ҥ�	yE�4�jp�r�X��j�D�Ě/qF��5e�я�Kd�ʕgʵ�O.�ⷓ0/u�d�)�d�����0�n�	�}t��8̟����O��m�z��I��J3N!C���EQ�X����^��.v���7����R*Ѥ�O��{O|=�]wq6���p(�D�[�������`q�TCٲ`�`�6��ʜ���o>�����=�B�jOe���e"%4N�C�i�Fu�\��R��F]�4��пkkn�rT�|��)PY'Z��A�5w���������1����A�dߧD�	�W�P&E�Ďs��z(��7kbDA}�gn�U���<O��1P�F�R�;@ͱyG8ع�LBA�N���.�5F�/hea�.\�-�$۲h��� �&�:,��z�����=������Q+���1�L}������oʭ��8����Zu8�g;�Vy|���Ʊ�I�l�7c	�l?��3�J��I1G��.�w�l��5�)����E��jiS"��I���B6m�M��7�r|Ώ	n
� o!W7b�_9��.��ix��M*��Z0�8�� �*�nHz���첳���De�m���%�3���ِ�JG��)��,Z;j������O�ٯ�
�w*՞U���:W�Wzc�$j��B�<�eF�Ue�Q�*�B�����s�.1{)G�޹��`  ��(e�$��)�T��ߦ�,G2�3?D��7QXf��D�EmL`
,D"!��u��.�<Ʊ�);�����L�aE���z�(Q�(Z`<bU9������*����+ π�.�F%���T'��Oe��4�,n@C���V,����8�
��G�S;	�?ù�'��r<� jb���yQ�q����32�Y21���FI��Ԝ��,g �|��-:Pk,M2	�'�.�J��X��*���Y9P^�ce8�
�I&
+$�R�-X�hA�	�a�o��L���l5��� {e,��%y �8����业��{�y���'�O�B���_�Bp�p�bU �	��qyM�� ^<κj��	�1ش�Q�bA���Z�ЋJ�`�x�[��(� P��&jfV� n}�;��/���#�n��]!��ʥ%�e�C�è��M�	[r؊�N��ل*�Ӑ�����]=F�$^u�����11� `H� +�P��^#uǳ�^oi�ԭ��wmg�j�w�Me	QO�{6Ђ�-��"M:t�ui�a1x�_[-_�s��0�����N�z	�]������9ܖxB~{�������`n4�l�ܪ8G�Ő�S6hx�ߏ��_o1�"4G�q�p�\�p�� ��=%A�oT�.@�R|��n_:� ]̹U���6aq栶�[��#��߁����aϪ��G+p8F:b�N5䠽�XTc���=	���xc�ohL�V�gؼ��E{(H��`��.=�lf���n?/̀f��G��G�� �D_vu�f�s!i������~F͖�O��H䇒�y�Q9���Hu ��!h/Ծ��)�ƙ�O����;��!�_�����p ��%M�����.]�xP�����3�{�]:��!�Wj�M�W@U�Rɇ#�Q�i�ֽO��a����l#PC�T�!*�N���&k�XR��� hL(G���[@|ֲ/m�����Y0l�Ϯ����ŧ�ºܝ��Gn�Z(J�Sc G�J�֧�pù�c��L�����C�*(��1ʟ���?��� ��#��k��V@l�&b3?�jP����+�PX}��LdEP_{�����4?�гs�:%_P�dRuy�"U�?���5k���"*3|k�c��FHv�]�V�e=�� @|�Ц��,���%H?]�O!�.��EX��ƺ�� BNÙ+�+��-"��Ғi���d�.A���c&����S��֬�/���滝V�1~�����K������^��d��*�fjU��/�y�޷�?�@�ۣ��ۖE`���c
3����+���I>����LK�}
(ihm|\�q��C��g^j�Q��˗Pht��YO�׿4��o�d^�����<7ZԐ�e��˜���F�+���kzdT����h#Qy�"$�6��Iq��b,=V�����uK}�+4���P���f:�r`֝bO�?��@�L�r�YC�7��U�@M���:�Z�V9���L�����)U]�,�`���F��X��'T�z���+��@=^�|о� (��2�<�z8�r����Y.���-�\�؊g�3P���f?�ٶe|v	h������Sț���;�3�{-Q�8?��th%��T�:�"O�U�ESr\���-Q�Y���}I �X��B�����i�9�a������|�Q޲��w�z�cU�� ��5�N����(���T�2g�9kM�9�\W$$5�E�B�s����`�AȾ���^�՛陷�}$��Z���b��n"�<��3�!œS�y$�d��4}��#hn�j	r)n���̀ߴS5J0���N����-��`�Z��'��σ��'��8 �=~]$��� O�őw�O��0z]��7�J�Y�����l��*��N[ysa�}�=w�RR�+CUL�sJ��az�m7�e��T#`���Sz>�&�v���N���� �FנrZ��#~υ��+�g��hɶSy��J�x�!��Y�#l|��ƈ$��b��	�C�W�Y��f�����K�Zf�2	���^�h��_ߖJ�#ZS�!5jQ�UA���X�T�	����*�^F�n�Xgƞa�U��@}x������U�iI���u���~I���� �y/mR�~�f��/U����r�]���l��9�f��5�����V���+��tW����W�(k�u��>dʣ���^�5h����՗E��)}4��k�J>������;�\U�m���jj{������Ъ~�+��qc���7�m�"�+W�g��Q�n�D������R��sY�FQ�ӛ�gA�M����F=��jo�c�ٲh��C��; �+��-��.)"�iq��ZU	b�@�K�+9�q�ף�����-KcOX�>ڶH�-�7R碅����ブ����=��?�Q�̸��=�*�����������
�^�ڤ^�駞e��Bhj��5��e9P�\�-:��/?�pI��,qwW�A�m-�^�5��'v�h/|��vA�v�+�~�-��
Q�2��܌eA�r_�s41���z���a�&&Ģ���Z���UX,k�M[5y#������C*>���v�7ï���-�ح(U���4�?5-�E�:�[W���ދ��o��#h!X��������M!�bUg,�;�ҥp���D{��1
�D���cGP��.
պ�?#)�3�S�q�����)4�T"�EdF_�(��p�U�^6�.C9H܌��D2|�����V�F�6��7ٵ��Wּ	�>����g� :% ��_μ�0�\>C@���d�J!�I%W�b��Խ{��P"�l����1+1������l*݆�����ݻN	op���!�-��l�H-����$3p����?�|º�o!�F�g)��(�T��b�a�pR��[�ӫ�CV83�P���yo��hEy9�G8cEn��zE�����l��z��J4����X�)�����_�f3tØ�NO�l�����2f�jQa�\ڼY�WQ�Q�ѐ:�ʅU�pi�0�1B_��`��4��@iP�&�t�b�=�,�X0id�̎7�|��̰d�@(���m��w�e�f�a
gM���ڡEI�c%2�'O_q��jBӯHu+3�ks�D}��*�o�  2��j�'+ O.ݖϷa[¬F�M�4g�$�[u��T<�<��3c���V�U��E����� ܞ 'V����-�;W��mz�/9&�;{)e�n�	0Λ�l�~tr�2��څ�^A�z��E0�C�K{Y{��3�!�n��6�Au	"���p�OG����Ҿ�L��K�0����q�c��y. Y��F`wK�e�̬$�W`t/�=��pxԗ�nܪ��)��PM�n@z�2�I����E��yX�;	o�$�1����v ��� r (V���6�gQ�DX.x�J�����;QW������r6�7�~��`��S��d�gb,��\<d)9!`��h�t�x��%���.=� �R0��𬌰`jAW��S~Hd���0�a2nКE}^>�_�Z�v���L��5Z�PRI�SA��7���zIﶊD�T���z0w\n�æ��w�8�D���`E�� Ȳ�5�\zZ\#���|��V�
�cI��6�W�G�j|sAoE�` �^��Rк�AC�eg1L����2�Ro�
3�c�]�AR4��%b�s'��z�ٜ���/�#�U>��L�yT�'��E�d��M#À�T�q���%�A�[�Z��V<h�L'�գxq�]�t���P@���I0�-Z������I
L��e��x��$�c�~W�Iq'R_3�˵�xN��^_z����)�J?�t���Y�:����^*e$�"�F���i���^8�,gM8죆��������+y���6�N�=��Bn�a�E�Ii���I���&6E݂����X k\��/KGש����T��F\*@ЏqS i"Uc�f��k�F�a��3�BU/�L����`���D���q9Ӣ���1�V&HW�ןΩ�˪Γ*�e<���-S��s��ir�IkH�I���L�B�%ﯻ����e�K�%�3(�� m�2cOb�si�I}d��9��Ü�o.�&�������ʋk�t0s���	
�\�<��*����pifб-%�2ug��U��c���`	�_5gL�?��6�ʇK7���H�L\C��SC]�RS$��3W��Ђn����d'l��YHi���a��[P��m�b�MAv�
K���}��s��M8�GuW��i�]۴�8�nⓣ͎�x�unE�o@Z����3F����.���Р�VjWR�Uj�����R���/~����F	�Ymhb9C
�;�LH�U�\�J��py)+����0�&4 E3��j��G��Fc1)�km�~ps:���i�����u/O�_���iǽ�9R�u�mԺ��,?8"\=�7�F$W���O�/[=���� �ڍ�'�Y�Q�fN���0pLE4yz���h?6oB<%��.���l���{��>��E��\��!4��;2�^�~/�//�[2�J�PN�`�hi�V�7�#.��pݼ]���^��ء�rк�BtPz��.ޑ���8+_��*��U"��RB�p��a��O��J��HK ��;I�|�Y�s��u��t���Si��D��q�3�����ˬ���O�ÉH-�lo��LX��e7-�<(n��S#��� Ed<t�B�	�U��G��1��b�ɋ���=�Q�ᯖI����=��j/w!�p��(\AyY̥����;�|�M@,6	��m�M����*q��q�T���(�T�ڴ��r�f���,+C���=�!�/��%8(�Tv�Q��������ZHE��n�r�1Hr �ML���|���d����ft�t�1��
Ɍ<1@�,��HK�ߊ(���`�:=��+t�7�	*'P�G� ����߳6h\jJ�E�a���<e�Db�Y�[~�_�̷���?O��N�%9U.�-r8��V�b$�O~ⵣy<UX�`x.ː"�UO��X��T��͌�N�~'.�����<�m<5�w���f���'e��U�ƣGq�C��#��H`U��gF���#� ̡�]"�g�y�D�.2櫮��=t��	�}**D�|Hr|�����p\Ռ���
�˟��'�Xn��1FL0�l@X5��,8�X�J��� �e��6�"sZ�T"�<�4!�#�5������i�E4@�B�m�*���0�o��ꓓ+z�[?Q���%z̆�?��dUΧ�����"��|��$`P���sD[���-��.������h��J��5L[����@+6������(�Ͼr%�Qw�*Vg���A-���$8�/[�IY߼׆�� ꆒ���@�{�9�C�pApd��>n
�����%v'�\z�!� ��l�T��M�n|D��� c����J�(����'`ڑd97�2]Jw9ڮf��/�	5��Nc(@|���E�� �r)h����=ط��G�����F��ZD� ��?.�}��� �Cc]�b��;Mlz��.Ӓ��m:��d���U�Edm: �Gd�d�H��<��H(�/��
��)#���D@�\!�L��:=���Y8���4WDd��%'��U�6�u�<L�`�7��#f=?��?�E:�P�Sq0��8d����#U�B�d��#�ʖb��=D�b��3W�Z�.���jj#fʛ_=l4�P�/�_7�D�E��;C���c�r��-����7�)�B���T��V��L y���|h9����	�.(��3U%�16,K�^qeP�kx��y������Y"��U>WW{��J�|�$r����n�K-��� � R�|�U`��,��G��L����@à3~��y)���=9H���t�Û�t��W�/�a6YB�&��Ϻ�%��/A�Ԗ�����4Y.�#l��I֞R�)s���MD%�m��t�aC:<W?�	��vW�Pu���&�n�>;@d1��vS?�{�k8&���`���8uv@�d:�%>�}��C">Q���m�z4�V$e�c�
�]����Pv��_��(XF���m�W�r�J|d6^3�
�	���N���^K���5���}l�4��!u5)P�vM�������K�g��7=!��N#�i��(T��W>L����'�O̩{d��C�|�/���\��t�$�u�F<�#Z䥞��6H˫�z�S�b����2b񿶭܂�嶎�Ѷ�է:� �	(�ƣ�����:H�au ��ץ�2e�)H��)h���Q�c����a1͝&���xcVR,m��^<�C0���)���w�������r��W��\R͗F
0%�4�S,�y�cO4_���`b�R[	f�lD���t�7-��qd��qZ^���~����G��<�-8��/>����fI&S9Q�ę�r����Tf6ރ�l��6&7��c�r��J��8D�\�VT�0������Yp]EV�\�	o�j�]�Vq�ﾏ��'��J�Os�3��"]LQIc?��&��j=#�{�[|�o��kе��͖��XN�F�jy�e� `�>��]���qw��	[����n�Iuآ�E��-2��֏!��KZ �&';Xy��R�!4�V�	LQ/҅��א�?�EɎ�N(hm&zɷ�`Ck��i��"��B�0�zC����)�����\��x�0��ɛ^�#�����H���ꈊ>%s��;����� $O-u'anh�9��vk��͘���
n�.�����ɝt'O������
��YѴ�`~��4K���W��6ȓWv��<�+ٓ�MP����b�J,#��C���8	VO<O��#����؃���xʚfpU���DD�Z�7����|���垏���0�4��pe=^���gԜ3J��!UG����w��us������j�C ��}�a�7,+���B���[�.��m0T��h+�l�R�>5JAgz��̱o�ҧ#6�T��-K�&�8D�[�a�iT�]��E�H0��\��ٴ(�����M�0Ա௯7В��{���4"9���� #O�Szq�Ii�Ϯ����D�r/�k�T����82����y���C���76`�#1M��^�ˀ'tÊ]�y���e��+/pl�-4����=4zkt���NU�Q?˂�Gx	��@��lOq��6'+!�R��#�����)�{v��{�(`�����A�V2r�H"g+㣬�n���i�� څJ�p��z�I"Z��^�ɶ�@�*�Pz�@\�
�)\TB�IRL2y������&�El��W]X�,�"��<Ÿ�ѫ�Bu���"�j\�)���d��T+X����o�6�1CɓF{����+��L���ָ��#/����Ҩ�L�����_=�<��+mz��_�/�b�����&n���^� Snj��|Δ8+b�	;3a�1��|�����L@m�,��'"4F�*k~�?5���"i�2Lelz��Y!��0�raR=��T,�]�t���z$)���l�$q;�.K'�a�*aE���e$�>���?=@�ݴ��F�r�Dj��f@W�~oI����˖(P��u�qsU���bf��0`���
�uc��h<9�Qc�����V�z��q��oP��M`��A͊B��um�X��@'��(����²t�o��� ��v�{\�М"�>gzE�䚋��6�8�ySE�ox���F��yS�L��RD�K�7:����X�X�Q�&߱^P��W��ieY�o����ш����'��D��� �Lː@�EX4缋�(p���K��	v.zu8�F�C�m�3���U��1�cu�$�Q>��V�y{��d��^����Հ��j�&`�zx#��^�|&��.>���*0�4�G����e�i��\�-�i<.%G�	o�I�4e��b.�-ң}�Q^��r���7�"�^��6��'
`������2�XC ����K�w���:'k�E���6����E>����F�ae�	l�P��t�&}�
�Z0���/���3V7��ã�P-�9<�\�F��g,�-ȡ�&
v�{�&A��π;�1sP��P>.�*?��@��c�H�/�"6�ٱ[C�Р@��R���öO���٩ �ڮ��/:[���M�G�[�n�Ǜ�A�6�X7G�I6�,��-m*�8��5n`b"j��S��Da[�i���J�SJ�_xS���7:㺹)����`=@��W5ְG��4��Zƹ	�K#���nm=�+�Q�����r@]9�Б���[O�����`�80T��3hC�h������gx�8�473���E?�a��!S]�l��ûch�p��Y��Vʡ��	*���dU3����j�ѧ)�24_VUd:V���z�E�
Շ��^�
y��0����8�@J��Dd����;���C�:pa$M�rHP=�c����*��s���dT$�� ��O!�$I:�� ���o7	Ũw��Z�����XG�f.�p�
����5j���|
� ���V�V����D�~��f:�s����FS0��Kċ�p���K��1�4��A��U�V���Eő�8rg���T�Y�-tM�H�8��{ʻ�u�W�XT�t����qot�~�jU��5��U�A�\��!tBZb |n"t(l�}"�3 �byi"zXj���4f ��N<!�R7���-lv(��_��~xu,ǘRԣ�eJb#���L��e��8��[V>P���@�c�����%"y�NŅ`�X�*_�p�[�x�{<�-$y�>��^H����aԺ�s�7��0��s��{�dW�ҟ'���L�T�.L:�C�d��2K�s]ɦ>q��c��u"8r��5T!õcS�4��.&�V��-T/8� �G�1�j-�
��uw�xj;�b*A�~oyG�Kl�[�Hx;@�ݖ��HVK�A@4��E6����1�ZV�\����P�-?{�n�RN� +9�n�ppk8�>�o����y��KV�7S/��i>T��O�K��1U���/�����[�۶Du{5<�aZ&5^Vy=�����:2��,SAN��ի��${rC�r��:�$���rh�*T�y��9�U�.e[���`��{��RT���V��&��	Q��۔GD��.;��~�N�n����+Ġ�SJ�>�|��F��:B7��܎!�,��qU�Kz��ws4qs`��+T%��Np+/���%}tŋL��k{�	m��o��`��Gwm���MR�x���HPm���a�`��Z��a�{5�?UaQ��Zniy��voCg^����{b؟d�z��I�;�Oc򍉢ɉ�h�"�$�j���V�3�Ft^|b<� �:�թ��:l1u�
��gzb_����-5_��G�	K՞	.���F+�o�p� C�Ғ���� ����p�1VT��XPu�I� �����}�>�	�@��!�wF�tq���#��y���:��)Ae�^穆����A-�<���p��,�j�i+�)��
BC�oH0���>]�-�0�g?W[0,(l�zjo�Z�u���|��R@��-�[t3���K�U[u���aK����b���.�ԛ6�?W.�SFӫ�\��%�\~�s9�ǔ�\�a���QIż�ݕ	���0Fj����Ack�7z���{"�9CkFH7g�o���%����zަ$O�hʅ�8�/>�.���K�`e�UG�.����t��혜��S�;�2����l��z�^��]	uU�̳�}�����C�A>�	���@��vv}w�o�[��V���'��5�ͱ]?�\�[���~�I-N��"�6)|ꑵ��t�lq���4\$����M��l�+���L}�O*��Ob���D9����7���5�GD�c����w��(4��\2�y�]���j��@,�:R���
�K������;�������Th��E�LT�.�'�,Ñ��wVAe�Y;fܓ���[��<:G%�Ϥ��yo-�}$��^S�qN�g]���IO�
�����g�kۊu�7�U��4�]��F
��3G���'pi	]�����W��u!�#����#�,�#�I��^�>d`w��H�7A����M��&��#e���v�'{4J�7��N�4|��V�G�u7�A��b���{/��y`	�S��<Ja��##Z�a��O�$r���WGva<�ѼA�Ϩ����`7&���X*{=�0N�����B 1�%C�%�\k���<T������y�D����&�޸q��%�z��*J��{vJ���<����Gje	z�������XG2_�er�ɡXLU���.��>b���V��/3��(������N�+<���Z����Wcl���*�C���wHy{u�����o� ���V셩�������P���J>:���(�K����3q��ƦErD�6��Q�_=��%����������U����v����Q��}�;? ؚ���W����2ayg��)�V�5�ӆ�"rÇ�P������������i�Y?�}�@Q$�͕��y������ ��G�F*)-~�v?a�bh&X���f�xI�F+�Q�T�h�E���^�zb����`�����͓yy��b�-=w�|$D��(,�5T�SR�~�tiH��A�Y�T3�d0�|J�vPJ��$�������QI��7����M{��.�ٴ�J�	7�c �hh:p�`�,o�&:&X��GzP���'Q�w2!u����Gv��x 3<�枯^O��c�����\p�Y��(f��T�������@R�� #�Q-#/�8�3;# y�6���£�M6���.ra�lA�t�-�&��о�J��<6��z!$=����L���A���P'�;4���6���3/ML�"�Zo��C�����Tȝ"���p��P�X�ވC��e��hE�����&3�~+��T�*�qC�eŇ��G�9C��S@ȁ���n|&��UP6w�@5���WװȘJ��ا�N:�7�������ʟ;�0�"QF�p�r�8���P,פ��,\�d'��p�7��M���Q!��E1�N�Q	��Y��٢��!oO�������I9A����o���o��\���bS+
������S+���7H��Bx��T��Qэ+*���6�v;�����m#E�:�������y2;��*!~UjI��,�3����l��R&���|�p�z����t�r���$���:�jX;�ŤR�U06_�ӣB��ݝ�9�N0B�j<��AJfL��{G<�\��k� �dZ��ό����w5�:�/앯?ߕK�d���)f�u�)�x��_��o�9ZAr���l��i��&	 �0Ip�d/)���U���Q�'�Tz<�<�u�7��h]�d?��	���$V���/�4���7o��~�<zC�Y�ֻ4�e-C餑U��c&� ?<�8�W����+��;�s��ע�����J;#�?�g\$U����Qt���j��W�,��ךnY�"��"�>W\�?'�%_sV���@�}��S]Q?�Pdj(���bQ~-`Fn4>4ݳJ���l�A	���]����4�j��yM�RK�E5toЌ;d�&��şڙߕ��$hP�y�.�M��0,*4������	��"�]-�	q��=a�K��<�����h��ńL_�V��޾�n%7��سv��T	���QD>�}�6y�k}�
��|UGZ���o��+�F��$�_Kh�M��슏�F�l�8� \u"(=�!闸��x>ՈakI�gEc�)��^q4���q�{p)})@�(͓3)K��E�v|v�F��� �
A?:D�8ԧ�D5:8���AfqW0Z;����brzpb�%�:�X6�N���}��jj����-��)�氽��H�Z=�M�F
�lR���p��灉���g�f6�Yqgq��Ew����)��LBNh�ǟ��@¼���r��%e��!�?$M���E�8zn a��3%��f�m�c��������{.�Yeρ8༝]���*	jD>}?-�Cc�=թ��U_BA����q�y�2�5���c̣(�c��i[�Ζ�d����x��㰁ɿ����j���@]1ɖe�C]�)��� m�`u�������
�h�B�&/;�����2���0��V�^��8Fn����W��bֺ����=�zo��th]V��>�?�|������Zo5���1�?
V�gP�X��"��
'c$�9k�g�c(��"�2�?�rN�Km4%i�*B��Wz�F	?�܍_�c�' ��P1���p�`l�#p��