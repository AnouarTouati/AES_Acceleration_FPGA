��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&q$�7s-u���Rf�_M�[n������6Gw������'�sLƅLÕ��V�pl�����7�5�Z�[���������������t��K�=�B�����Qbx{�� ���E"1��,�`�����0����bOe����������-N���X���v�W.����h�o-G�蔧�tS�'��`n6�����f7,��8����J6|X��� ��=���� �Qbig��ɒ��-�z�j�'ګ�_�(��ޤ�qp遼�<�e��L�mܫg3����~]sR���yF�KƟhYR�cFb���V;̸�{`G|~���?��@ȶ�Y�P��xթh�ꈊ'���v�M��4��)�,��"�2���xS���`�0��㺽ɪ�L���Y�O�ᑈԎh~%�V)[�~~��U�FBa��uc�H�Du��z��UG���!@D�����-qj/�n�V!�U�z>E�G��H+:,���@�G�����mcyH'���bu���&��h���˽�JJf�~^�胇E`�\��8��P>�����>��wʟk`�)%����Q"��QN%�
����c�z)�����ז��pZ��!Pawת��9�K<N�Zڧ��4+�a��}4�P���Z4[G�{���X�jX��h^����#g�䉿��{�ۓO��Bd�MK߰�'=���L�Mqu��(AJN?OH�)la�o�6����ݨ(];/bm�C#�-[���M؇@WX�f0���(���0�?��K��q�+�41M�>�(����Ա����\R}@
���\�욘2���\3��p��%l#��]Ot|�X#g�0�Ən�aL�#�¹3n��Z$W���\��G��)�904ևF����˵د��
�x��R?��.o*�����A�S�W,�~���m��(XT���V{s�?fc�:$�xމ��V�X���;Ҡ��ta�N/�΂���Ŗ-��B}ɺ&ӷ�� ����y)3r�3���65�\�PS���ۡ�9�o. �d��&��M�#Io�N��y��7PV8s�-���V�5��
|�wIq��\�S�W�o�O�oT$�(O���!⡄�+4	�T0l�&��cmW��V�%�.�&s@�WMq�S�z3vP[?�aq@��+�OW��Q(آ���Iޫ<��S��<�i�����j��.6j��K
�X�D�$��W�xU:���w(��Ő?���Ch�pm-aw�@�}��g�q�d����FeB&������/_��&������9@1��Z��"է
4c �[�G1l/9�j�*D�l���m2,�+ K��y*T�9�q�ّΝ]V�B9C�LF�|O3��l��3��e(�ʨ��E�W�YϡOĴ��Z5��`D�����^��EW�M{�Vz��6�����t��/���_�j/�=C"�w��y��r�H|S����Cn�dҶ�b���Tp�}��#��C�!ԀXރ��|�,�vP���:�n\ l�t�2�`��?Y�-v ����Tw��;�wF<�+�!�� f��F��%�g���/��J`Z���h{�|��*Dh�K�>P����B.���Yvp�{���������_�0��&��y�����>ﰞQ� ��	�\����.ͮ��Թ��Z��Y:d���<ah_�΁ah�-M�-����]%A9�y�?�P�ˎ�0Di��ty��Z?s!Q<�^+x=˺ �kX����0�L�S��K�8�0���;����;f���E���Z�:���N˛����Y�~l+M� R�F�s�ڐֺ@�p�ͥ�a���~aF�T �"�8R��^����d>kΰ�B��K\���uN��>e���#c�'`����iP�a����x�B�\�f:��J!=@�� g��(A,�Q	f\z��!���96{���Z�xS��Y���:��d��Y�=�.\ݸ|q����VؚDL �V!�[04��sW)�54��rz.Q����/�ʙݚ��;�P��=ԕo{ ���g�@qx��b��)P~���D��^��F2�� wc�z��[��'n]c�Oձ�:��gA�4�o��B&������UVׅ�FoZk��z
�E��i�,��ǔ���&Tv.:E�d�i�D��`�uA|	���SD�>��:yi�+n,)<g_���w�{�X>Ǜ�F��kL�η�����>�3���+�� pz��rh�uZ��� {�y���U�"��W��S�Q���Yڋ�Bd�D(���fC��J|H���_T�R��������I�<>�-s+ƚ$35j�
�5-u�w}.�� ����(4*<5c|�+	���#��g�[q��+�/�W!��=h�{���������FK�f̥�]��a.�[�n��z��q$ECMʌ8q�翞��]Q�!R�y`y[�M���l%t�^�y�+}  �@��hį)%PH ���E���P<[Dd�TiJ��%�><f��O"���iD��tY�/�H�|���)ln��ʐ��Uu�#V�e����z������)3��|hK\�J�!R�=4@�W�"�`Oj�g�2Rl
�4OŇ~�a��:*��>wq�-��ч>�ſ���<ř�d�@ �-����G��O��������3A6���j���6}*�P�h�w`��/{4��3)�gQ*xʧ8*u���
����p_�Xg*cT���Z�?�����ļ�����)�-C�*	� z'F�!A�� f��L�><��^���q1�����ѭ�jr�.y}�iX�y�Ry��%�;Bo��\���6��ŧ.�i�X~\��1�'ec*Kl��U2�b�ق�F����ҏ~zk���9�=����<A@⎆�=���C�g����J�"܌QvR�Z]6�c���ֶ3a�G ��x��V/����E5<߳�m ߐ4�k؅;�%�V.�g��\ ��yhM�5V΋f��4���`g,t\\ J7�VR�#D&��Q�rV�L)�?�D��@��Fm
�s�ᲈ؃q��l:�}�3��y��~���,}�o�����$azH
��x2'r���Ώ�����H�ի�Lý���P@��FI �oU)��k��17�D�L�12�&;�9�U�[4�$CF�Ҕ�3�c25�(L�v�c0�V�2ϲb`����� Ƹ�ľX��D�6ް�p�(���۪�sK�[�6y�4ސt�W7�.�"JS���|&�}�&�Y�
W�ˏ>ȭf��.e&�-d�j�\�)�1�
�"�OS�V~i��)�G�1�Ƙ&0ǀ������k��m̀j��}=��϶d���F�e7�u������;�Fd&M���&�����U������Y��Z�;x/Y�P��OD��"����t�j��C#6�ǋ�����y��u!䲭tP�񂅹�N�Wk�T�(qXG߹�7���+���0ס7�R� 9�w���O��Ts��tMﯬ|%�U�9�^���:�J�R�ڇc�*��K��-ni/c���PeBI�W}?e��A���&�}8��-���(b�`�m�	����$�S�O���8w)����܄�)��D�<@6�#�
�R���|j҃����(�L��'�C?0C��g�!|e�1q�S���#1�2���|�$0�o@=d�?e��ɶ	+�s߿Px�h��E��%v}g����M݆N���g U�5�NSB�lC�����	<Xٝamr�*���*v�����]N���L�E��S�~�S�핗����7�h���%E�S����6k���ڝ�:�usXK��C�P�)��P�ZDs�<Lm|�$��A���P��������E�d�8�:I��K)1�> ��@m[YI
�4�&��yYO-�e�$�Ǒ�5�\�v����i�`O�%�|�o���ƚ�:ð�"w4ӶS� �zप����֙�c�y�"p,����*�8p��	0�lX� �2-]f:u{�U�2u�os��P w7p7�H��t�����?7s�3{*&p�Q��7�HVo���3��3A�X�B��쟅[a��t�Z� �R �kwQ�͍��Cvp�}~>�j4�?.�~��-mSQK�.&��I@��_���6,���M��W��$8���,: cg�iS�*$�`��ϊmhX<�k��<�E/څ��,8gP�R![�U�~�p���lT����$e2K, :a���o����x��G�iD"v=�j�S�&� ��퓓��Y��s�2
�3(���/w�i�l|���l%��$t�^ji�U΍�G�_><D��b�;Kqs�`
u)���/=�;��y�sp�<܅fd1b&��GK�<[�G�M���
UQl| v�y/
���{H6M=��~L/.�m�	�m�Wo� �R��Iu%ܫ��t���g���d)���>�.L���$����9�j�V�G��w� +�Wޒ�*���	���K�=S���ĔvT���z@E�cf=]
IV0"�ͧ�V��$������Bi@>�.���g�h	=�Y�C*f�q��r��S[�֖-ܑ{e%�MK̷<�}�%ȩ� ��[�C�:���+��:<��bxs���\X������ĵ�D); b��v��'�l|ïm��G��03h(��f�Do�̷Y}Ӻ&�h�h��	J<*�|��i��pj_�i�^��Hlʘ&��x��[���E���,���xV��1׊�5�^&�Z�!g^�� .D-���%#z:B6�R�M�n�_ǒ�s����D�x�DS�������Pj���*�9��3����+�������޽(�V����G����̩���M�_�F�~*HжR������M���x�b�l�PL���#�7�yW2zg@�ggw{#:����h ���ݙl�.��֤�����N�vp�ڍӮV������y����C2*̟�w9��Ahw��𷽜G�H;ضUY.Ei�:�K��W��o"���/bf
�uG�	4��]�U�������Ée�i�k��7#�8O�	da;�c�]���%T�P˾k*v�'���� ׾Ϫ�y#� AN�М��6�|�<��$)
�x�Ԕ�Q��״u.ᚌ#��G���� ���K0�w�� ��M�r�=қI,�pn��QZ��6/s�㯞�*ꢠ�m|�2�\� N/�Yx].`�(�b������J��{�7ؑ�6��6�	:U[�8\Z�)����[=c�P�^�%p��}h"�]s�.�p�
"���8墎0����wބt8~��SW��8��{;ږX{,b���tF^6�-�n�V�;g����>Y�>�$���B������������ŵj2�I�rybk�(ə�`[�0A���9%�΁@D�7��5 ��o�����B;5�uZ-�����}��WѼ��u� ��h���`0�# �Nrf?�YIA�Y]��͟�
qA�3��E$�f��tv�/\�@��*g~��VwJ���*6%�9U�5׋o�W+�q��#�W�Yrl޻�\e��^<� �l
��:��R*��<2�]�M3[x�k�]v��K|
��VzE"�{��+M�Q
�_�`�1|��]+�Y�7����Ad���W^�b���_'C��d]I�1�%e_mi��ܑ�"Tu iY�>���l��HcQ��2Oɡ���%a�l���]��~!������t�!�j�  ��k�Dd'}�[�9(&ɫJ��Э+f��oƝ�u`�N�aD���B����.
�XKTp.��7vp)��8 �v8��j�,e���[|�ґ0�Ïڨt���X��:��l�>y ��'��y�a�����4��?��]��븛�8=�1�.��Soz3ܼ�"��e_�/�B�������:��{�Ajh����'m`���cCm��Z��{��|�P�gq��!��G.���%����e�Ç.�i.l�9�'3�N�/��acޫI:���ǾB���~�����3U��I]��*]��}��S�ꭖ�U�����AD7��$�����j��l��Fw�*�meT�|������³���^ݍ�>����By�a�r����0��1����^o��O��qi�G~0�a�K�>� �<c����m���V�SA
#��]�<n�/9݉�xye�AUu��+�������M\g���e����*����~��.�H�n���YB�y���u�"J:��IDuqV	��yyy<�\�B�T�\��\�K��¤�橫����"��V"=�Y��n����H͂z*���\۪<05[g[�����</m�iS0��f:(�
��h.�Î�!��\~���YfN� ��1�9,�� x�E�d~ ����z+T�(�X�c���D�V�"�h��\��*�4f,P('B�D�ܱ����-��<C��f��B�Ρe;|���n~���@�dA������Έ��I�)��D�R��.��`��}1��c}��b���na�Uc&�Yl0cX[�
�(�L�fp�E��'7��w�O?�(�B�w>?>z���@Υ�����@Lg�:+�
L{Fg�(��Z��aq䖤s���!�d���ڥ�b �:���%\����wLw�H5L���➏7�v=�6唕�B��EɌ����\��������#o�R����H���e�u6�[7�>���r?s�����.((��p��RI3Ĝǂ�$$�%8���_�+V�`�-�[#���W�#}@z���ήs�r�rM#���7J�n�^��O%�xU�&ȝM�[5,����=C'�QV�ʄ�@��
�ߕ���o�M`�!o�|Y�����M�Jԩo�o���������3V�6��F��_@��g��V�;������C�u�$��+6�}���`��k{Yk����o��cT��A�	�dW)b5>�NCт����M��N�RZ0���D����%I�.����f�i�#��&��X�#����V�{�]_D����+�ٹq��C�*Jnה�B�GG0j�`���h���!���ô���SRv�I��U���m�?)>X\Ե����k����m�Do��V ��'�YZ�?��9�IuO۟;�z��+oG�^���R9Z�T�e�X C�h�l
��f�!m��]^_p��5~#Tʎ5��st{��+�0Q���5���,X��	rDN�?|����YC�c��SbC;���|qޅlj�ȫ>s[���h��n���^��;4�p����$ҿ`wr(���v�VTe����b��k�;	�k����V%�6�+-`�kS��1��i�u�U��8g"N?(����7��o�Q]#{�+�m�jk=J�!�x�P�[IaX��T���g��e���6�kf�$`�U��_�����Bf�/������*�-�yOJn�=�h�}���@� Q~�ii�л3�<��t�'�6�{�lFf`P#	���H���1��� ��Q��G��W@�m�Hq^��-�
����Sh��ӱ��	g�^T��bY[��i��N�Is�j��a����3�}_O�6f�۪��S�_��O���. ��S/��klv���N�iN��}�I��g���M|<�m&ڲ�T�C�
���yF���8���P	Z�������J�4�(eq�P�j�k9,)B�i
3��B^�
`��y��vI�,h�6�d��l�6���["�يe<Z(_<p#����TCv���i���;�~s�%.K"���%����*�t1����!e��05>K�Vq��0��md{��a?p���Sh	�������-��������|��>9�#��ઘ7�|m�zr����6��G�@�A����۫$>},�F��ގi@ȡ��e��<u�v�9�f�\�U)Q���Y����'����7{�+��7ꩊ� A�v|VZT/�]��b�s��l#�
T���0�rD_<kL�B�|a���V7��ҕ�8�]����c�)ﹼ�dQ�_K��C�h��c��۟�<K8Y��$���"�f7<�t�B�4����Ձ�����v�B5��:�������;��d��j(���Ŵ"�p���Vh�G-����ZE�x4a��7J���Ѧ��{�e2�3"L��r����I�-�t��/ǉ���GP�L�@�图Bz�n�`M|�2�қ1���?����_uU����-�������n�Ɋ;\�%��eJ�WLh7��$�!</�0�
Õ�dE�${-i	+�������X�p%�7��5�}<wQV5���~���E��a%l��C���C�P ����ظ��b�ͮ�
36b2֕��Yc�D��*~X���|&{q��wFzG�ȄL�p^�!�N�+��:L`��Z�������'G����Zj�~�Ǣi����:�Em�yP��Zy���yo�������� �Q����m��d
5hX?ܒ
d#�.]7@+��E�.�*��$���x
k"�}zJU=5Dr��r�ZƼ*�;���e9eR���r[���ؔq?����<�;/�ͻ(�Ro@���b���i�'��!�0���O�s8�]1+�=����')|��ֽ[⁘���.��H[T�\�!����1(TԎT�H��ˈI&Q:��^}�F��y�OF��~��˕�4!v<q��|)�֩ҿf$�?w���!�,�&H�l��{ ��O� ��%���d�Y&ճ�q��^��(�b����W�B�ཌྷ<g��و�8��l�Bg��Y\��po�ba͢E�r�-�҆0j�4�x��J4�O��/�Y � �q�u
y�{�4�v���^mlcx��Äh�^GO��|���������v��zē&�r|z��a�,.#�hd�����q
we6���1����1U���<�qg��B����2U��Im��3�R�^)���1�;b�ܞ`�v�4V���Ϲ��@P�EBLNr��	�KG�!>ל�̑�Ⴆ�ԓ�7�v��*�qJI��3�������dT�aa�����d&0q�`kEݙ�;�9b�����_r��9V+7a�]�m7!���&΅��Q��e�|ۧ�|�#���n��`�=��ó	/}i�1��(���y�5`���vr��!�33:���b�eL����P�
��~��"	G:�4AɃ}:���)��֪'��@-ැ�~��	7R�(q#P��2B��Yd�1�^Ћv�m��3����X����IU" EB��c�Y�=S޼����/��P~�F��dY	�d�?(��%� zn!a-{SW��I�E��A�=�
��"��b}��!j�Fm>9�#6j���u�9!Fx�Ce�1l�N�@��%_K���U21�8��L�����.�$�8��K��E$hU�<����?,�|�j�\0���/A��;&Kt�9�2�5v�߱���G�0��f�ϊyn`@܎b��y���駵����6O)y��}�z��E�ꖹ��H2��,"'Ux�b�,��ѷ:Y2��c�|sc��_V���%o<˳x�bCU�q�,��+���Ǩ�(��/���	^ұ��销Ro��I+ƍ��\�lR<A���gG��@\a�PCg�7k
��_��.�o��L�������D�}�؊8����S�Uy�8J���1is�e��c8 >3���~�n��3�^���⢜aX,�ۂ�N&���h�Ue<w�G�������R�
�^GMR �
z,M�=��D1Y�'��a�n<�<K���,?�f�n<B?_�q��:
"�h`Q��3��Ck�k�'�S_M!�aq��X�:��"Q���v���'���<\��O���>K�u���yf���w֍��%b��8^w�Z�@җ�{�s �z�d-��eo�R[�s5�2�q�X��<mwb;�t��Yek�y�T��Y��9��NM��Jev��Qh���dAС:��4ߍ6���R);�x=�}����~{���G-�֪mc*��%�tw����*@�C�
O$zW��z���!g���J&����e��.������O�y���s���gXq���R��������"Z ��E�N��9�:������H ��/w5�є�%g���c��E�MU�~����i�����sLC@?u�,���Ve ��5�=�&v��_�M���+�?��èA�u� ����w��J���j�<�V<v-� ��ҫ b���` 4��U���F=E�>A�9S$�{�==Ɗ[)����I�Rbނ�$�>�#���iSb�8�WB����qCh,�<�����#����� ��(/4z�8 �+����7	Z��h��c�18�A�wY~�1��J��Fp������0D �Jv��#��}�r;�eu�^)�'�>�p�����Q	;�ٗ�C֔���,���<'�,a�^�k��}jR���!�+�������4Je��mo�N�H���0ڽ���w��y
��4*�����^��6�8�o��|xȒH�*�0����ѵ�f�'C�a�?�ch:k;lf��g^�Wx"��W]lӰ��^��h6h�+�J��"��o����y�n�+��_?�BN]7��C?E�9XO+}��o;�د\���T��[6esam�S�����5��s"_k�e�
��1���¯� �t]�?��Rg�]=$b������"�L�Q�|E>H���ˏ@U�;<�s�#hgm����Ɲ��D�"dtD�rEX�������>�7!���̱�!����A���7��LL�-��]5Pt�ni+��1U�lu�k�B�T�ζ�-1�%�eثiu�ö_��i�g�2�NH��]����8́\:�M���xbpq��h���fD櫓2���l(L��hg��g�X?�}`��<խ-Wd�_���E���xb����}� ḽ1�aN�Mp��ߒ�,�J�_!#n��X�:�`^vU<��(O�NkԼ�~�!�3��7"�ts`y��l@g��BgV�Q�j_��DM��e�}�!tJ�������:��H�u{��{2�F$�k��6�\p�-,�\�,32[Q���6m�v`H��}UO0F9(d!��Z�5) G�-��C���~U���v�[�}�kb"�>��T�����ֵM��Zg,yt`h�6���	n,L�6\P��y�k��C���LA��)�Uz:-=H�␁6��G�����;#N8�)�L�G�Ng4�]>���ǕM�����oFjb)�<�i�B��Z��W ���~�d�B@W��fr��(H��c�2�C!�) ]�B��ZNu�jk- �`
��ڙ[e#�7T8[��N�="���* !���G%Y��:#g�y����.�G�s�ABT��[�%�|[�y�$�IG�g�@�ӿ c�qҏ���;bhv^��8���A��]6����=�K~���蔴m�����SM�.A�pS�*NRYA�_���}�?��m,F�;9�Fz"(3�R�b��dЮ�
�{U�j2���`�����=I�,>���Fux��^�vy�m�慆�Z˾��r��v��6Ah���|ZN�h�	��k�S�bpѥCTekc��+�)�>6��&R� ��J�CF��k�䍺{ɬ�z*"�n
��v��X}�o��,����Jm�u����iTZj������`��:�Ƒ�zJ�Dw[ԝ�����ES˓f	�f��!��waf���Z>о:�r���j�ދm�ñ�"��2G�b@���� J@�B]���#�#ms�,�s(�*H0��g@���w��1
�ZC�GG�dX� ��Kݗ���$��`C%��Z�b��@1��vL�$b�|�k�'�"6�ZV�Z�|˝fH([u,w9��94��-Xz;�VȚZ��l����[���d��=��I�d+����]��Q���)������i4>{��I\�ݹ^b%,@�p���e�u��E�;;:�ۘjs{��� ����Kvt�\�y������{�'�!*7������Eq����������춊���=I����"w$�	�γ	nG|�c���(5&b<��Hb�_���ai@�+*A�_�?�8(t1�Y���b9���Ԣ=\�n�<�|����b�w|���}Ӊ.K��b��j5�Zn�e\�*��Ò��P���\_A�-�	�W��cy[I�q��m� '��L� ��$�����~�C>�٣+R��7��5b�L�k�U�mg0|W�/�ŕY�[��<4)��dW7\.��LZ�+(a�b\���G<��(��y� �4,��]X ����)�������x�_��ߝ=i�*��#7��_��Ėn�e�%�GY6E�u襸*!m�*4�^�,�<b�!���}�{�����she#���'�ֽ��ȧ�����X��+ �he���^���k�¨ݽ�bm&�h����Ʌ�~P�+E�davz@&LCJc_!�y٢��]����a