��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&Ű��=�b��vT6�4��fWg)l]��@��7�B݂Dۉ�{��m"ԴT��L]Ε1���ɩ�����B���_��m�5���8��z�ߩt.��]FNH���V��u���|�i�$��#hHR�+�W�lN�m�ǌ�A��ݰB4��z����(���Ec�d���+v��|���oT�ĩ�P�n@[4���Jf����c�V�o�`� ���Iޱ���h4 � 9
Nq+�Z�'7t��p�-Xp.����SY@p-s���*K�(��� *$����r�#̤�:� }��	����R<d��\@7b���0^P���9�p �� �n�]���T��� 
8�X5��
ι=&Z��m?�<��j~`Ñ��6�+(��W��L^bW�c�� ���-:�b?�B�8F�y�R��/�?�Н�`	v]ҹ��ҁ��j
ӡH�7A*���d����Ui5ku�*�E֢}�J$'�0�Ś��$PlƐ�=��[�%C�)J�-��Q�S)Yoȷ��Z��#�V\��	Viz�k*F����".���DCK>X�K��̖�ݢS�03�̿g_�T�;c%��ζ9�N�)����v���-��z��.R��Vwz���{���ڌ��C�<t[Dh;��j�;9 E��j�xO=S7�%�`	�ms�V��{~>����{�l�5��^M(,e�rss����#���ĕ�H���L�Ǆ�����e�h�8d�@	�I:X�iCL>����2b�](����*�R�,�m���0b�	-��ړDÑǌE�Vhn�����E~pϺߐB�r�|Yn�<�i�?�˪R�z�7�RO�ۦK6T	8�3�3T&ߛ�U/���+�&X�j�Tؗ���ׂ0�^A�s�܆�%)!ل�:�}��$e| cp����0�B� J`��9~�Y=��y�cp��_;����&
���Φé�����TO7{���Ж�!e(�Ӕ��"T����w��<���S��A��ڏ�wf�@}�gy��H..��I%��D��<1���8ȟc�� �H���4$�؄�}�u�Xm5��%[�d�m��C	��'V����\"��s�n�J�@6��߳��{���!L{���N�`%^����9�c,f���
���K$ft�=v&ؐ�bb�#���h���	�n�xT]� �\w�AD������'�$I�,[�O;ф��UOj���'vo3�e�t��F�cy�/�����J����QU�ƽ~����� t��蘠���t�����Mdf&�����Aq��h�E�%��	�U����lc�a�I.�0��>��N|Ms"(U+�+X��Fܨ��<��wr�C>7g)kyG�}xw�m
w���ѕ�X�$�?�,}���+�b�T��Ȝ]S]O��0��'��Q�4y�l1ٟ~�rڰn����.�V�̕�Z1	N����V��4�CB?��L�>$N.�V���F8,a�/j���f�o�+l$���WW�td�G�h�H����:�D+�]���!�@��Z�7/*[��̕��|��9z�;��5�(>W�=�M�iY�SEP�sZ��^�8�D��;�_��L)�.��!�(�B�׻� Y��7樓���'ԃݗq�$�v��Ǒ�t�6W��S�3[cW~eD���$#<�֨�RXPh�j�3xɹ,�� B�@�% ���p���{~��0_tll��x��pI#�[�c�bxﻘ d�,pT8��M��׫��6K��N��H�k�@g�������Sed���ۘ�v\��̻���Gbuz!
�ぶ��߳_��TU�VZ��w$`��PDßrA5�u{T�t�܄���~�E��%��E!�P���z�jSĄ�_@�GD���>d��	]2ٍl�3���n�
�1�;<$"Ua�'��`�I���S��ba*�vO���za�rmN[r���~��I=�{72�K��?.����U�ޥ"&��Y�TD�G�tč�އ�7��k) 4�l��v%�u�r��J�B4`�s���J{�����|�ӝ{�K��:U}���L�c;@�ԣ���O/��{ɨ$=�|����I5�c`Ӳ�`*nǿ��s	�Ѐ����v;nq��8��PMx&����Z�BO�Q��y��X7����G�-AQR�C!bϥ譋�p�)��J�!�]/LI�7]eB�� �f�S+87Fd�ECv �#��tت�C���oIh�� �NR+��L!���Z�B�(����C(������R�J����Ա��|���8���q���h��XV��Μ� ?D��#���1Vn�vW��,���\ï&+��&gf����|\�,-�ɸJUڢ}��6�2%�<�ms�a7����;���F��nvH5L�cZ����A]��*���=&�);�5��ܾ�aq-��̔2k����]	�bZ%�_{n/Nُ�(��ɋF9��;��t�?-,�6�uw�
q���f���%�At�й9.N|<,�uг��<�<�EƲ2����FqOw�˿���G�Xi��\��C_A*��,ݟ�a �w�n��@+%Lއ�$�Ms�WY>��`r�Kd��4S'���d���=U���G�����:q<��?ё��Y$��N��Vo�tȱa�%-C��;��c��wtY�	V<[�4����}޹u��mC���O7�K?�\OP�By�V�C2͓����u5�������LW\~n�Wb׺���������gҽt�D'��X<A��1aw���Ł��M���	��_r�n~)�@��#W��z:�����Χ�Q�Nq�_|�"�"l�kԀ����>7dЎ��y��fX��˸;x]��>r-1��+�e�fҲ}�d���	��.+�e��N$�s�ob��?��	�=�W���&6�t��B�>�Ff�@�bvb�꾧{�٩D�*��Ә�i:��i�>�����y��8��ֆ4��4���Ni~�~��f,#�aE�"��N����}�7�:Ϳ��og��U�(Xsr��$m�|7V�z,r���G��
ω����A8�ac����$�+�&W��Ud����{�I��4u�;��TB�l�ۙ�y<dwl�!�	��i�ܲa3en�c$���o�m���ǒ��G4[��g�^�xˊ!~�;� ��j��Ҷ5�MsZ@o��Re(��?�Z���A�-��"�⮊fۡ&٨t1a[��2K�s��t+}g૽f��ݦ���DMo���=��X+�Q�{���ECq|�~��G1�SBWM���d܀.��ːQk!�1}�n�j�E!''��K�AwJ$�k.������f�3�oO��%��(��7}-
���"+�~긪���`�%�I��RT�����_8*I��5�0�NZɷH}�)NaŸ�i����9)�1Nd��Щ�ؙq����P��v�q�˰/���)�
S��D���ye�tEc[P<8>��[�~�X~ N<[u1�V��<�|q��-����`(���k�`�O�f�-��l�l��@�-lβ3����c�,��@[������"�a�̾}̨M}��X0�V��Eת�$�;9+�GH#@Qz����L��%soc�u�V�l�u"��'i>��\��@<gmM�*�@��p^3dU �,�쫈�����, x�vϬ=���7�ٙ�Qz��h��!D3�#nj�j���Fc���(�i�8\��QV�u�X��3~���^����l����y#+����.�o#lV��Kx��`��vD�R�z1k�ɚæC{��>��z�!�e�z�T 3���Ib#~1�dݠ�����C^#͟�P���d�@�go�x�N�/IC�Nr�Ѻ�<E �ŨS`Br�7E���A�9;������mN�o�qR}ӯ}o�ӟ������J�㖣�E�5�?���JC�>�]֠�B����|�b,�K��Y���S�ζk����9��H�Q�JGH��z����R����p��Ϛ}-|[A���!}�Nzۦ�����B��Ǉ�.W1�|N�%��I}u2P�1*)hr����B�Hjͥ��>���jz�l`4����
��)<�Z�.#
�Wrɟ�)7#@�x�E�L�6��\k*N�c-���}�t��]d*].a��[s�>����ty�u�>�H}).q�V?9�'-5!�9�K�L����v]�M��[R���߷�[E�f&�;p3 ��p�Ow�G1���*'���<̺
�HG��y��v��].p������W�:��S�O+y�x�=�xˣ��9��PC�*ˡ�LHDr�p�Eu8�"�_�yr��	{����6�o�c�(%ճGa��Kk�@����76\:����ў�1��|'$�N���0�7��9�R�5CoN��@�}֜�%�3�3`��d���zWw)���[.��z��n��8�aCՍ��	N`�e`���^0���@L��}nF�����t�g[u�:��:I��A���ԁs'j�[>/�AƱ�[6?�~�ڊX(�Kmf��0s'�a���IT��ޮ��T��>��w�mQ��FB��[9b[0��Ks�^������4��R��ē�a4adH��$��	���eբ���I���y-s@c�d����~�9�$�p���L�h?�i�os���w	_��ZJ�������oH��GոVd�2�9�jq9���I���U��,����m�H��3��I���[@�r�ʎ>���a�R�!�G-��R}G�?��*f�����/Kp�t*.���F^1�Bv!`}��ע����%�����9���U���2H`Z�C\�?/bZ��y���Y=̈SzC�4�W���M�]-L'������ �y���;K�qx����Z=S�!�����T��`�@7�t��?po�����M���C���՚3�8-��0��P�Gf��zw�GH�o�8��@�*���~:\��"��.Od��4]��%7C�d%y9X	��X��R~�s"l�d�K��L�R�zs��ާ�4�i~y "�l��Y��B�[���o>WPd��9�
��A��/{�����#���ۿO�g��A,3E�i�����< �k+�̿U������o��t��	Vɬ>/��I�	6�����|)�}��V�����oQ���u��e�7t��"�Y|�ڂ�DxY� ������_��z6�p�_Uʭ��xS����NjoLT��ן��O����� ��re�}�H��ʜ�?e�%j��\�/�0����/PL�]��):��e�o=i�R4�O��p�1#b��K��in�g�N���v'_L�*���,�l��N��y)�ǝ�����a@~���Q�R
�a�8�򙒏�1&�(5������Ovd%X�����ו�Fp�^%1��I⹣*�������;�@�ݸ��)���|}h�*�%#�lh����`/����!hpXh�`Ȁ	Ön~�;l���}���7ˬd���#02�g����K�Nm�� �D939�>�q`��p�b;tS�X;�y(N@��vtYv�:�CE��Omm��� ��짃��|pY�����RD��W�	9�J��u���sPX����H*�b���O$T[�ag6���,/�&�<��ک\�9K�ɩ`9�U��F����L�� ���}I�����0W�����?B��{��7u����\S��8F�N^�������D~����x�լd�̅6��kѐ>�Ykx#� ��p�R��ܠ~��3���oǎax,f��=���
��'S��\T���y�]�����Z/M}����U�h��޺�|nf4W��i�Y����\q�y(g�Ps�������
O���|u�v������ѓ��RPL7�\��Xr}}�P�M�b�%�W�!a9���(z����zu,y;�KF��p��(�_CU�I=i�[�R��t8�ʟʇ�(��Q��6���Z{�A���M��V��4Իaӣ���滅��%l0B�bD�Cᖱf%�+�/1�E;�e"e��A�T���#N�|D�>�Ao���|`_Ƣ����8]��Bv�J.N��\A{F?1p��cU���������ړ܇�P�ԜSȐQ��@����}�:7^�ÖqD�B�jFZ�Gx���]���59!�'�?�A��ʢȳ����v�"}S����7��kYq��c�
d���s}��Z@!g�p�<��@A-+莩ka�U4V�:��)%�bw{�ʛ�I`�K0ۥ�d[������T�.�u�
 ?�����$���WX+�a����(��n;��6K�З
�x�G,^��	5�n[�ƭ��\�Η[����I:��gקG$�Z�q�R�rXuT��6�x{+��|�f�扈�eTĵ<�^�2-��I���Hf���u�m���"��=0w��~���d��6j$�>B���K������"��sې�����_�cX��Q�rD�S��L�ױQ�:8!�[��	Bg������!��ƻ�l��jW+�b6-_&r!/��<kW�+8�+v��kcKb��������^:���=�8<ߜ>���D��^�wsX�^Lq�x �E3�}<��Y�29�<�yE:�*I���Q2�`,�
.�Vp�(Q}ME��,�ړ�Em�U�1jE�u�Te��14��=:
��4���ISG`��l���3p�D��f��L��n�>w�еF݌�q�<�`>U"E��^�F*ʺv�?�?�����P�[<��%`B��#FOM�8ͬ�*%���RϴX�#�f��uE@{b
�Rk_��[���[j�Ҥ� �s�ӣ�5��M;�rsz��۱��"���)�O�-�����U�t�;����
��<�h'�ݙ�ӳ�����b�}����?�Q^�%A�[��
1�~R~7�L���(�v�)nA�v� ��A+f*�}��8\ �R�p.-컅�!�
pV���cJ0�EJ����Bh�-�"��^��uW�e'�_�	��0ۮ����9�~�р\��^ei7иDZk�+�$Ԧ��`�Wc,�f�J�Մ��Ob�����c����T�٭Y�Q��X�&�O�t��j�x	����������c� &٣���}���Q�����W;�}��в�0:�K���d�����6x��J%�//9|��];�^���]=A���F��N�IʫO������o�E.f�������������Y_`���-l%V�v&޺�"-*��E��e�l	��q�p&uu�k�A��Y�
y�*���Bگ(PJ��z��#��K[�jk8N:v���3�N $���싁ޭ�L���ϋ�S�E��K�v8P�.���ۛ�uD��D�^p[$F��ZQ_LXNs�f��Ew�o���ET�4��{P�i[ C�D���U۵�;�ziT�O̽!r�����*�>�=�,'��b4�vWWiM��1.�r��r�h�����~D{�+��Gq>Ů��<ꩂ���m{1d��d��0O�����5%]�#�𮟜�#@�0���{=}��&g��=����R�zA�����xv�kne<I�m������Ӷ���)%���\���{����hT.pa�%kߺ�a�|_T5�O꩎�T�=��#�i	g(e�����7���-z
��`^�_��N4�)k<e�J���"a����ɩ�j��2����d�ߦڟ�Q�5�?��GR�(+I��)7��YO���f�u�L���/*�B5�yG`ٹ��%K"��H���z��6�]} 2�qfxć�,J{,�aGT�	��yd���o�AWeã���Eh��?P�A T��?	�9K$��n^��T#����0"�,oX�S' ò��Z2u��ե^<��w�#&<ڬ��0ʔ��H����V<h�ï�����+y���'�˘�'xͿS��Iu�Rx�Ox��6J]w S��8���+���ޒ�,�l��<	6�z33�q�����M�F@vA��p:3_l��-��êf� i�������+Un�k���l�{
b���yt�� B�����}�k��^�z��U��T�m~%֐�@�W�
�&ID>�|_��6�Y�St�N��']����4W�c"��s~ц�M�X���?J��H�Fh*�<�����3����%�&h���~ǝa�zDM�#��隑��������n�/|���-�i<���� o�l�-�^��D)�a�f�������d�xtaa}��Xj������T>/<1���pקrD�x�0\���ơ�oD�&!l @�ߐ�ed��*���G����X�ږ�D 50�
R 4�jH.H� �s�@'�y�v%^T�ѽ�H\��2*�����>�IW�sH���4��  �Urg�_O ���q��,�M:!�����5(a�_̂�g1R�]L+�ϣ����En�j��9��P�Fe�wu�Y�tX�N�"�*l@�y���@s� t�q ݨ�𙲄U�P{���=����"ts^W'"R�\�0��?{�^ ���J~�)y�}}�� �s����9��-�����[��j�xæ�ȉ]&0g+RM��=��4ǭ��~���E"��H&B.���!q=;҂� ����.�#��T�9�`��kIt}?:��N��9��Ei��2�����.��޲tK��o�ܩ�֙�?�Fz��'/+�ӑ�;ϝ��kC� ����H}8ʡ���|5
 ��f�e�<��#��>����2N��ʩ ^^2�X��W�.Fg��fR��3����o�Zb�d�h�h��\&��,ℊ��x����W�`�`8҆��E�w�ջm�G�V���i�ڇ��\�)�,8VNxa�~hr*گm�fi��qX!��@��=�`���������:R�$d��/թ�����;�����
�t����F�z��Q��s;�����������Ҫ$�ClBIjG'��y�ըbi�[eF�q`���F�&]���x��oM=KY����Q�"g�;��xq�踶����3�ku;@00���']N�V\�[=�0�o��6DVє��s���B�N�8ڲ�T���}��&9�<$�V-��{�֧'6 rF���яJ. ���=:J�Q"����^ӱT�?�U�Ե&֐#��>2��h�zm)lT[���r+�#������^���5��y�K	{�w��jw���D�S�3T��kc�=1�3��R{(.�sf�t�Y�c�@��G~A����TA,.!@sO�@U6^3ra,Ƙ�(�R��5#tl�y�������0�9.t�>#�6[�ܬX�G�j΂�� ʠ�*��.�x_���WN*1��,H�+�u%�+g�dǫ� �#y�WBt����ֹz�F���
��'f&M�w����$:_.����6{㼔�tCڻ�O�5�ⰵ�Ի�3���w���|�D�zd�[�����J�9Et|>�*�:v�Q�\J�_?#t��Y.ۼ'<7,dd����J)a��07H ���n˞=��a�h{AD ��@��!�a���>[��^�sxz)Ra��<���W��neL����GBp�է�����i��M�*�D65��'3�-� U�@��g7�
@�G�z*�X�Mig���Ⱦ3C�G}��!����%9(V��W��U�Iv���N�\C�7Ґu�B}?�݆P��շ"
�����$B	��O�F���� 6��5L'�|�.��Δ�z�j�[�o�܁�_P�ei���ݺ�_%w����@�)\�s���V�ac�6�jIN�P&�[1�8�1p�A�Na�>o9_��)i�f��'M�#�f>�z�.�$l����A��M����L����&�����zwB�	�@�;x�Eefa�#�I`�m#��kB`*%@���3���D^	1 !��/�D�)�f���Ǜ�Z��%bQ}9�g�����l�2e�����2�T�ۅpo�o0�_��������۞�0�p�<��q^��p�bh�d�{Zi~�M���'�/-���/�� ��#��Ϳ��5����7ח��L��71&��v��i@�U,"������@H�@���I��E��cZ�ʷ�،昕F�F��z�����R����p���ǒ���Z	�%���C��X��R����Q�nll�'�� �=�ex�FPV�������n�ҡ �Q��%zn�F��a��dtQ0��Jd���<�	NUg�Ĥݛ�S��3%��Ij���Ӓ��I Z`���}����,'s�@~`�,@�����oYi��U��J��5Z����I�^��\W]��݀��!7T�b�=�-c:f�(�48F�j>^��/co
zj?����ݱ��*"��>��2�؇���G����*���Ȼ1��Qf�)S��O7�o�.i$C!5��.���5�|I����^�el��l���	f�ơ����twu/p���R��%楫�����Ӆ]�6��3ET��4�Ё�:E�mX��~��AX��ڰ�����TmA�!���0��Lu����WC�[j�E�uM�F3������,��)K-��/��@�3Lv��kB"U-5��s�m�/si�N߆: ��7���'8qyj	��g9�M�l!G��Z�t)4�5���xy��?�mV�����dݲ^�,q�<�z�q��2�+VT�i�܏���X9*�;�a?�ߠn]�Ș��k��ǈ~1�'�C��~^��GfY�u��6moz����9;��x���gLz���osM�H��~ʠ(
�0������Qxqq�b5NG#bMa�*�Zp ]N����_��j��am�Ҏ�r�7'��0�~TNCҌ�5ܘ���l�1��\5�ܑJah�ziIßr���\>H-�������3���S���`p�UZ�Q��3�^v��d�z'�m�B�'�����)i	��k��c��o "-=%zIi�[������]p�n	U�ЋI�L���1z��F~�W8�Z�M��N�m���(�̿�o�q����}��	���2F�V|�AM�\�� n���J���7C}�;�ܹ��KC 8�Ɯ�CYR���.VIa���+c��!���RT�C��C��.QF��	 �D_�6.%�ԓiy���R@����L=�ow�;U%�3����<��<h��G(X����%1�r�H=X-�����a��nHv�&sf��a�g�urN�,7=���z�ēC��H���y7~��<�O��-D�8�UXո���p��݃.�[���͕��h���.��Ato�P������G��o�j,�gk�e��EdV�Z�Y�@�p��ư�>�����v�*�-�Fo�0S>'���Z>�'{�4�5m�%9��j����I�"(j�Q�4�z�667��g(��7�b�~�����Yň�:��*����_�/���AG�Fs��A��X튀��#yt��#�~�b��
b�w=ª�	��\���ƶ��C�hʋ߁-)���ߑ*]�r9�a�P7��l_MT��[~B�*�Y۴�&3҅��|{Q���O�x��%���(�('[J����˔��S�B&�X��ч	>*~��r�^���G�-5 �<�ah��f=�ܲ*��*S�\��n%��!+*�b�P���$0��m�_	�e[����e*��&����m�e-,��i�G�K��
�� �:B ZN������3�`����p�3����3�c���]�&Ѽ"�R%L��ĹY/^~@;u�wi<�,AU6���U����������oV�h�����T4|��7���zt�D��x������|���	��C��}�=+QB#����r[{�x\���w�tO8Zt"R�����2$=f��6�=-5�q�y� o�2�2x\���l�8�:
h^�|�h�#5�U�m=��cb����rw{{ekr+f��u�v�f�k	 �0C���]]}�{�����d�w��칮��3��4�@>a��k���HJ F#��|`I(�u�K�F*�8������Ǌ��rҠ(�k�Wc�p�����!8)	s�V�������,��,�	J��.vl�'?�l)�7�|Z�l\�B�dS4��%ο�k���Ì���<���Hv5K�� �}�]t;Ė�{�?##��3�5�t�'��y�'�jQ�.����twp��O܁~����bYoe"�М���fp�{Z���A��i����P
��e �`fI�[U|d�^s�-fc���F2�Ȫ�2_T��=m��캅�,f��K[iWR$��"�<?ab3@z6��y�D�d
����oc�D�Q�tb�!}�M���Q�����1�-M��2�x�e�_���ƭ�_����L��~W��1�r[Yp�q*�"�d�yL0�8���"Z��J�	my����XBTB����xJ�W��
@���SG���s����t��0�i�A�<�,H��m���k���ػ����A/�\i�[���X�����S��|\�՛��c�&�m�YU���T��?�f&T��1q+ԙ��9�]2�r�yb�X��R���+�yq��t0� �=r�����Ն�U�éP�j�Y5��������;(~t����?�$Ǥ�A�O�w���i�,�� ޳i�_�pgn�y�����$���Gxj�3��+c)x׫��Qx�)�Y�M�κ��u���QH��fw�ėN>f(����B�޹뽸.�m����G?e��u�e	�n�ˌ�>C�-7Nś\���	=k�Q4�Fg�:v���A�D�Ѽ/�B�&}h�6i���$��w�
���U������9'��T���67�?�`�[�Ts����y�b��y�,�E5�`ש�H�1������R��wA��B�g�4�<��1�
��<�pk�Z$|ͤ����L�ϯ����G�4� !�ܶ�6q]�alXA������<�R�C� %h�����M|.�E̛;:�[w�=WC��Q
P�"���
^"J��0�=2���bPK��������x��ĥ�(�g!*ޏ�o����6O��ğ�PD�2��ݝ��@��V�Pԩ����|Bb
��@�s�%ędA޼,�i:��l���$QQߴ����Ϙ^mⱻ��X!��7�����4����H� G
[lY���d�n�����j/���F]ߐC˻�Y��(�M<͒U+-�z�L�o����v<6��z��9-�68��6�1�H��H���Y);�5� b��t�P��z�m�K<Wb$ h�m���\݌U�ϕ��GG���~v"=ܖ~��L�%��̑��m�b��*�aP�䫱<N��$� cr��4���d?�[� �;mK���c��&$Q4��Խq�bT:�b�ϡ�sq�3Ƕ�׫?u����'m�3���*5�B����:��p:w�x�.��l*`���lc<�8�i	�ai�;�d���ۑ�)��%cgF�#��2�p6\������I����	ي�@��� z��"��9�lO�X��-�7b�y�?��|(e�c)>����0Շ�N0@F��d����\� �zF�Bg��E�Ď޽g�Ӥ�FUN�,,���}��٥`�p�
e@�T�iS�$ ����Y����m�`�u�b�|� �����ۤ��aS df�%��˹oF��?�Bk_=��9��U)=�G�Vi�����%U�>O���ؐ���E�������fMs�(��cU���z�n�s���@.O"� �FӖ@X$��W&�j�^�gO@Dm؉!{��W�R_Wvm�S� ��:�1[�3����a'�*��U�d���f؅�9�J��j4dt痠
��~"� �v�boP�@\�F1��r̢v=Ql#6�b�v4�\Δ���~�<���FPT3R�y�X��a��o?� U�ʈ���x:
��l�#�Z{@C|��9���G��v 
NW��:>Ks��i�j�(���{�.3�hl	l-^������}W�UfŞ�����dx��]��fʉ�g�ጟ�/$�q
v���e��������R�����H>��tW3�3�Wˋ!3�a+�a�U#�`7GS �u�uʭ��ۤk�C v���K������1s7\ޘ;Si(��YؖNF4M��1φ�����}&^}`4��}WHl�C�ǋ'��%US������@D�h*n� E&�h*�fV���X�}����i��l�L/�jE����	�]���4*!e���,ymӉ�=������ߕ�/+2@��rà	j�QsL��+�����0��ؘ�%tN��)]�:�������Q79����{̟��۸��ȁ��0y�`N[�;���e��a��n�)D��F��\�d�����`���h�G��W�K;38ݥ�Fw�E��+h�����J�T3m��kߙ�z!�PHB��h[��r]Xު`-55���Wlu��N	�J*~7fց�t$ޠMv&��SFh�#�pN��v�}e���g4ˁ��2qՊ�5�Y�/��;��h$��hS /QP��H�J��slD�X���'�&eE��\K��:��p�����ӭ�
7�u�R5��7���FԏѪ#�b�O�o&�l��0��A]��[���/��V#��]��{3�-3�?+�L��ˏ�^z��ߢ]�dt�h'3���?a�7����Sm�~�,���d�W���X���J��.~a�/�̢!���%�9M��@��ѯ���Cl-���Uo��
JL���I'�J~y��|+=����΢�6��a*�?����D����Bg>� �j���M��&�_[���F�R���ᾐ͵�0�^R9�T2��p�|��r!����ۄ@j߼��Q��oXO0nW���v�>�L��0A��-s� y4����S@!���0��B6��-"��A-�}d HЩJ�»���ڑ��Y������Q���h��{{�o�^���|��ׯ0��x��à垡���b#'�iǰn�"�=N���!���r9Vv�k&��DS�ӌ�5!=�	p��F��!DQ���S!�yf^>�;��J��P�<���G�V7�2ne{�9c�?K|��6µ�O�z�+G�Q����}V��	8���3�2w�?Ɩk!+�ϔ[�ǩ#�f"g)������Q������_"$D�=L,�#�����?��:!��.�Jl]E��mk���vAL��V�8`G2	��,W��(�k�q�%��������p�>z������/�z}�0�c�wk�w��(�3q�������Rn�똘t�>��>3{��U5Q�.&��e�u���Ů	�B@���	�`<:R�'Py�p$ֈ���˰nA;�KI%�ހn=�)�wB�}U�~a:؂�";��H�=����^y�ʹN�Ѿ��!�r�/5ki:X�%J��Y�LEMW���+��Q���-�8}b|�����Sd3@m[c:��E]�J�O�j��eוC#����6g���se):�s�	�[���$x�H�\Rnݠ���O�D�N�z�A�'lㄆP\G�i+˰�ц����Lo3h|G�&�2�1D	���u��'�Y����QTO������s��F}������%�>+�E�x������5��N�g���y5ޙ%����
Dj�&���-bЦWW�&i�~�۶�$��ǡ,gX�PW.��wɬ�jl6��M��_c��-��n}����[m.ȫE���������p4�=~�����U'�3���wI�6x�<�)��m;�o)���%Y���op�x#ʘ���,iF�
CHc���<�b�t��i��u��wjm�G���P�7�B�rGK��O��K:�K�:���na|e��؏���)�~�:�.D�O�����с^v:K=�/%���F�i�:\:;����.ڧ�4fo�+�<S�5����5����('�ГX��:+��Y��E=���h�D?o�ǽC.���i��I��
㫫�M'em�3%k��˗�	/�ި܍M�i2�t:�d��	!���9#���t̥��9
&��^�q�F}�n��~F��#�@��]Qٯ�W2�P��嵤�+��_���	D�a�סU����_|4\K.��Tv�_�v�W(��G,��<�E�&+����`��dE�Cz�����O�n���}l�����_��u�٦\��I�>�g?���`z�퀮�������7ܝD���n��{$ch���������s�F���)��lh�L��ʜ���@K��Lʔ9�_�E��|�N���X��2g60L%ɇ#u��)��j�Ȃ�WYz�R-����[��+���"�����D��,-P��d��������	V���m�����|>(�,��p���D@o�&��M|���sOro��|�4b�P����cQ�(x2�T���{�6�3�����A��v�X��r��pԗ��d�"x|2��;r��W����R�sҚ�JM��7E�,;���<gR_+�) �LV�lt,L�HUo��"7�&2�5�֊�l��fW�G�d��/&PX������e�������v��ҋ�|�M�ߌ�+.Ɏb�.4Y�0LH*3G���~�M�/:��7�׬h��	���LSvR�"ּg�G�A,RK�@������"����(V.G�k���ʌr�P�(�,y8��@Zй��`i"�e�#�dh�_���ESt���U\����b��M�ݬ1��I�q� RQN�v��rI�*��>�$��
q@��
��zS"���t���Pad��R�Č�7?�"H~��+����K&�&��hϡ� K�Qd���5��&-e�����>@���K���5�� �%���m뷊���d���C6�K��=M�C�`��ڽ�k����z�h�)A� ��n�X��u�d�~j�+��A}AqL�-c0J��qi�Cm�\�7�|*Gү�Q��e���G�A��v_>�	� �_�ֳ���)��z,��h�:#�3��� [�D��p��pV��&�8Β��&#hjӶ�AF���^�}���۲�x6�H��);
�����x�'��u�������e�pZ\�&�ֻ��W��8aK	��ѹs�bd�Ơ�ǯ]x�U����|�zR�z{�I$�K�g��lDt��;���S���'���.*�Z��DӍ^
�cxJ6R�R�٢��r0
G��(񍭓��7&��v���n.�!��])����*�q�J��4�W{���z�,�!%iKڑЦȴ/�3��_���!qt���Ҍ��zlpڅ�P��LG6��:/���_�k;)�p0 ���n��ą���*��\�{��xOH5��1�&�ʫ�y����}}�{2�Ƒ����*$�M���P1%)2���dU(l�O����|�U��к4�c��uQЪ]�C����tm�1*[i@+*�\υ���l�4�"®`I�Ń*rA���iSy���(}``^`�@Y����/�������_�B�>�G�1�h�S����d��3�J ���Η?��G��'.�Mz
I	�ң���`)��}��r�4b����%y���~#.4/z��2&�a0�c�g'|WeFQ~�G(�ɾz��{�+,i��!�����ܭ)^p��&�ѵ��U�R�)���e0[�U4s�������[ş��jd��7���a��r�y�./��،2�@!d&��d�,��H� �(�mm�pUk���g����e֔Tz(�J�L�>�m��������.2Q���%W�M#c�����5��XZ6`��Ϸ��)�ԏ����-Q��Hg�D	T�g���ג�;��$�E�j.#7�a�X� ���\~=ыV?��\D��wWH�SD����Қ�ZC����8/��E��b�s���u���7�&��ЙD#񨳲�E$f�d��@>�~��ȿ��ɔ2�HTX�"����Ĥ�����y({��3x������2v�!���X)���#,Af��V(� �}�(�S��%���,�u�W�4v���O�jTZ����y�޾ d��XNx���;=�Uu�ᚼ�hA�鍭#7���.����R���ڣT��Y1��Y9����3z��ML�a�"�������8'^��V�e�ђ͑7��:{m��-hd *��fb3i+C&�%��Mn묁�tjp�xKO�b���%��?S��1?�jd�%RR��6�l�1�����7�wzO��?��!��H,i�h	A��	TӺw*6NȾ���Q�u�|����!���A{ uEm(��xD@��\��r8sb֧��s]�2�6$[��,�xK@��
h�A�E��mDzn7��"ڰ��f��6qcՕRP�oIK�T�F�}T�Ί�\W��u:{���Vkw�|�L%��(��F�Urx�1���`	%jƫ�9�q_�sH�{h,S�_;�`봫���lnY�vۀ����l/��V${�Y6�\x�nXP8���w�� !����j��Қ39 ��Ƭ�q sB�W�"����H�D��xYr��2�oX�0��w(ݕ%:�f:O�~@b�7&����n�@Kݢ�׸����S���8�t�A�{�R�p�����V`��!D�6��H{�Q��5D<14�Ӡ� �T>���}�R�
j����8�I�:�yt`?R~��#�#-�JK�_�,�݉R{�<�����=��s�F:�Z�l� �y�f���I��'�b�B������or��0:�͹iު!���Wp�3ɡy��$B�T\���}�����r�v9��3U3:e��H��_)���U8A
]��l���eM���o��W�Z����n��,��X)���̎x�ߺ%o�>�\�Zn�^�Z�~��9�Hgg�b�I��C�p�C��'��qLM�G���i��{~�;������=lT6��R�\��1'6#�1��E�)ù��s�_(�
ڑ!Gw�H��c���U��hu�ɞ�������S0m��L^���-Q�3����T(ϰ�����%��;�6�a��WoG<0:*,W<�	�w?��L��LeK�����L�j�G�V���=~^}�U<���M��9���7P��9��m�r�Xߨ�T�l����
�}
%ݮ9݆����A����z�UnQ��l��hhL����}��N��V����%q����IN�4$3��M���]��u_-�f�O��7�U��Ր���Mǳ��:�Z���}�«�u/	�oe�U��8�7�ޙ|9������yT�z~P����$ f�\�C�ZN2=�I	��?�+1 ���&
�*�����%���9by���Gĥ٨�Σͯ.��o�i��;�>1�)���/�z3�L��E4n�E0�.
 ^O4���v�Yuw��g�f �̧��;N���I��<�@^�ñ��=��7�޶O�#�� 
��V'�,�h��Z�)���,v\�7��m*���9<�h�G��N\Q^����jy�q���h"��&/q�T��ʾ �iP�1�+�ӧ�����/0�zcQ�!w�0'G}E�_��k=�.st*#l嗛���������X5W:�A[ bN�)���g$'�B�1�p����0qZ�1�!%�M��e����ۋ�A��P5=�ܣ@����G�1 vU*m��u	��J&��a�(��v�2�����!�P/,�T}*�<���į7,&�u�^����{���q?sa�G�5���ݕW�Q���_�͈I��cV��kŪzط�=u`�ޣyoL�.���洙���uu�w_�Z���y�Su�v�����<1s�iЙ�SJ.����u�o#T�G���|m��A~A;<��#Ѓ�<�e��N�x�w!u��F0��?WP���ٓB}d�E����>DU�@�ī/�]�đ��m�ތ\Ǯ��u~����F��d�f�ɤm���ZN��Ƃ��lv$�P��w���/+c �����`t2���*�õj>&ݓ&G������*��[�i+]�2X�s�W�5��d/��3Ihb��ڄ���2>�6QZ�����Waʓ�
��G���6��ӏK��y,-��/��UdP����y� �˸0�%؏}�VH#��w��	����� W����_Su��
1z5���c��k�1�����]�/�ti���xن�y�	C<���*��,�OK\z���3�Q <���eB�'��
�ʓ�c5�錺iG$���I��W7�+���T(g&��+��Z4����=2����.�D�R���(]�&l4q�y�����oԦ�o��/��\Pl���fZ3zZ�`'���1��m�GB�GE�LeK��u7�X�ؓ�$r~2G�~&��H|���?�l���8B{�%�◦�%ְ`T$b�e������rAx�����Jz�Oބ���FJ�rM��=X9�t����s�l��(�L�T����$�-���B}��y���= �~�,�ڍ�K�g�Xp[�R�@��	1��%9o��ʏ� >OE��Q�_�2�\��x�ӭ�f�S$�֪ㆪ�N�I܎K�b�B�~����գQ�̼��[0��"�����F�ve�Y�$Ǭ�����s��ը�C�Ԩ�R���Y��Y�B�w��t�y;R��~��#�Mw?�<(E�<��5��/.�ѥC=�h/�Շ]����G>ȯ8��	��y����D��@	�x��l�ӓW�FZC�Zr��|Q*��}Tr&��p�Th�,"�I"R���ꌭ�]��@��U#�=�R�jv�L�Fy2WڎC�k\-�1f����OM�<Az�ߩ��aT�1B���"t�b���Ԉ�mm:��s�b�g�^C�� å��.ĉ%�ʌ$�ͥM�a3�\���k��	tz~�Cx-�P��'T{d�&q��劺џԲ��4�b��IQ��HmC�r�~��,wT}�yY]�����.�$��4��-#��j�)��W(Ϣ~��*�eX*u5	Ke2�B�z�1u�g��.���:�r�L��Ju�0�N7�!�R�M5���J����=��Մ����c���L����1+T*G�D��MqҠC�r���NM�R_R""�:�c9$ܪ���.�t�ʦ��b�x�f7fפ�ؓ豹��l߬�,�'���>��s�T�6���� �@�b���'����oV2'l��G��vRw�����+fg�U"�Y�?=<9Mq�a���s�qa�'�9Յo�lA�2��t���ᔭ����;���7R�ʩ�)࠳%ju��i�u-6n-J�/�^��^l���v����̬�jmLt� '�6-��:עB��/��T^}�t��HQ��0��ޥiA�QV���-�>R�\��*�^a ��8\��)�]��w&W�q�;�ŷmV��:�^*���4lc3&T�B��X'ź%7{@�X�
�0=|e�ԔD��fy')0�efߣ\�� vѣa��\i �V*hs��|��cDn���n��R1�h'���ӕt倒	 mL�-�d<��P ,<�M�}͟���b{emrmW@J���u�2�׷�f!ߡ�
����%4).K�}�� X�tLy M�$�{����@*�b�p᝔�RBك�4I�8KZ��jD�CN��F�K���oS)ۦ�b࡞��N���=s\�6�t�~��9�����9�Y%z\Mƺt���R
���g9�@�k	N�PP��Xz2Ey��rn�bL͜?Ҧ�<�1�	�;GIʴ2���3)i�|L��*���f�~�IeV��׆���-`kN1�U�����Ď�/G�eD�h�U�z�)�C\"��}AS8��+
��N$1�丝��+��GQI��_���ӊ��w�6ĥ�7�y\�,�;ih�i�u��DZ���_	��-���!�f����K�e3�dL��V��#����J2EA���Ի�k���~����A���^�7��� �HX'#��S��d��d�>)��Mfȿ�c�.J��uAa���������Y�W��F�cW��l2 ��-��p��૜M[�E�t����x����J�/��K���#�T_�����!���� �vz�6�S©k;oZ��0^�玙�z�5Q�$'p��.gn���w���ou`�$�]Y�h���5�*�r�0>�������K�ş���(d	��2�T]����Y����ey����:8-[��2���(4y+@�$d Zgh�_Il]�r1��T+����D.b[���؄;�>��S}��( p�>zS`�e�sF���㶃��%���}��$��綕���^�O�%���Ą.x�M�Q��K]*���e?��է3&<�mjA��d��PA�|�uZ}��ʰ0m�������L�Q&��"�xJc����d�қO���Sg���~���(�3��|=
��L�Tg��Q��p+'�Y�)+�S�F��J�T\������s��[��Zl�rE�O�+;�ş���u[+Xf&�o?M�H�R�R�"WN˶�ě�=>�V"��fp}��X��m����(�1����Uq�N��PW ��|�&��W�ҭ�3P(����L���]�3*h�T�<H(���fh�(x�F�>I ɫ�I�T�ζ�n�+�6L3�'i�_EP�Il�e/��A�[�h;9�j�'�f�$�_�J:���=w�Z����%�(��Ofl�� ?e���;�O��D�u�����\�	�:O��酁�k�� �e��7�#O����d���r�ȫ��n�?�6��u�l7Økn���;X6~u�����1*�h o��t��ں��'�6UQ;��"&}Z	�$��r���փ�q��q6qC�hI8�+���Z�RYڟ�Ї��"�i6l=t~�-;β6L�&����j��q���l�V��=�kj������RD��˞�t����Z�A��zJ1`�܄U2��ֺ�~�a�W=�����n���4]��`��:*~PI��o
}|�=*�����$Xa��O+9���F�>�D�0�HOo�Տ=NR�&Ķ1Bo���zK�x�w��s�{A@��f���[�� �I�"��2�m)�y�?ۄh�W=^�j�igI�3��=Tx�9M��Vy55���m��{G��h� �xƞƆ��*9�O�!H8���	�z�~�'ߖńu�4M�Q����U�Sx�c	D?ȫ�.!�F記؞x��yQ��3�u��u7��Ȏ��� ����^��q�Ї�l���`�V3�+�u�1 QMx(k��ՓNܛv�OJH�(T�+�5��p?ս�y4�lO!��[�RN�5n8��&٨��T�F���N���QA�^ ��ȣ��3K8V���|�b0gÇ��d0�= %x��k<�Z��$��J�o@�Bꗦ����M�u���)1�����7��a�G��&�)T�c��c�����,�_�GHɇ�I�D���NLt� ���y�l�Y����{"9'���WE���A5���at��u1�>$EpZ/lr)7һ��E�.׌ry�i&�L�p���b%����� c��x�-�q�C'�$�P<z�:��,�qax݊*���'�#e5�r	O��E�{������Y�ч-^G�$A�Y	C�C�5��Q<XW��/������Kx�1��ϝ�o�<����ߤ��ӉAg��v�Z�@1b�X���z�!�f2��mv=�">��C!�2�<���<�m��A�Lu�.�����Q�L����G�m��SS<�P�F偃�sgg5���9���A5s����Lfȯ��I�5ܡøb{Ω ��E�N��Z��fi���)����x���ҶN�DX'��X��T�o1˲�mI��(��s
�͈�'��m�v�
eiTu��[cjUH��WE������u҂��}�&��6����K��f}C�Z k����PcX�1x{�%Ĩ��`:��Y��RWI9̔!��^l��Mb��نB�T1����/ ���<�w)�6ٜ@42dx���3Rͱ:
��Ur�f(�1���c��W9PN�<�<"HF��Pu�8�G�ٴ��R�������	�7l'��A��HQ����kM0�� ��g�/���0�e5�u�,|bP=���k�<�~J��y-Q{��f�e���a��r~��T2��G������.q���u��ʡ�ۧ��M�z��Vjf�$�k�e������RB<�;/�NZ�c����n�4���� �\��@C���±N��9��a�;g�O�/�4m��������<܍�����������Z��૥\w��8��\ɲ$5�]�V��v�5��~ʒGx���%��9���*�~��t@��fսci�_`���2�Nw8���.I�ߑkY9�� #ٖqkm�f5k(d�O���{���n��|\-O���?Pl􂘭�.(�F����Gj��{�1�V�|�qt[�W&�"^׈��	����TV羮~�]U��:Fպ�N'U��;D,��S�w�:U�^�����Z�^x�g�,�e;�.���Q�lN��Vc�2\ջq�����:�)���
΃x��|ʕ�z�����y�}C��J�^�l�3o��YH����&������_<��%�ɦQuʎ�oZ뀶'T�,���/_כ7>�����������^D�2�� �8xK�h����2K�ϡ���rv
��e���y0`B
1�|�f	�ٌ9P����}6�*��`����T9Y�I�%�@�F��7Reoj�D�N�a�~"A2V ���{���d�̀�2�Y�"d|JE3&��?�>Z��@#Ŵ}�g����R�����{<��e���q�|ڧ97�5�)N����s {v>E�n.'��/c,��,[ڔ䷍�p8�亡�i6P����Y��A|v�����
�`���͘��c�Rb����J����h"_1��*���4>�O���m���Y9��7����JJ��	6yy��%2J�8Ȗu��PUj۔4�W�ל9��,K[A��Vo;���\5��B�w�w,e^wfq��U����K�.B�uk���Z��3��o;r���Kj(������\�H�Q*�s��k.�R&f�ߝ�ma�*�K-�w�d�D��We�#����b��9k ��;S)=���_{�W�/�4"|M*�*ʖ0���	�M�TJaP��C��� څ��!�,��8�x���Q9�[�'��U��]��m9r��u�?\[���fH9ԭc��HB����P��[v��f1��d��,����&�U���At�4��͋��s�5���w�T/&m��|h����J��ĳ�J���̊SA�p8�Q��ڱ3�n�ų���a1q������2�YdH�d^��7$�|����~�͐Iaq����*�����x���i�����OG���|�ɏT���S><�SR��������7=�Y���k6T&��o�؎�W�PίĽƣ:�����1��E��K�0w��} �����H[tn�
��"��Q��5�����h��?I�u�xZ0�)16���O��{��)q�q�gp����aR����iΧ썮l���{Wj:5+Z��j�2)[���`��?o<�Y\�⥴��0�����4�ƒP�T�����
�oMm*ܭ���n���o�z�;�#ϛ#QK�lcL��wޣx@ϐ���OMaWFҍ��� �CtN��!��"�u�5
�G��L�E��T�Xq��VG�mt��-��9�,6��)P�`�������y�Z�K�z�/k����yă�V���C�Y�s���Z\V��(�e�Ny/Ҭ��Z�R�����B�P'^��\$��ymT���y�Mu"�(�Ъו�m���*+E�h�e�",�v��+{����|ђ�c7��\W6/ߦqm��R�T@�1%�q������p ��:�a0�1��!G�.El��9l-%>���1T��t���
	�>�7�s�GcUs��^oj�*
C����{Ә�a�Q�Q�@rg[��,����_��Bk;�����>�ddv� ����j�\���To���-�ߙuX$i<�$��z�N�^8Q}�V�,`�8�gh��n�9sf8	לlt]z_�5� �"��zd�A�%����I���X��bx�����5u��j, D�9����͒||�J�D��J�-N�5���.>����P�x
�Xz@w6{�ѷ1�]\�mI�;n���X�
#�L�}r��YJLZ�kL�י��|t4	��d�5���.��7��p+�g�G �a��.�I&���9��,`b�&\%��ob���tm�
?f*?fz���&��eOP�sΝc��eF9���9��g�]O� `��&�������.9���u��yw�k��)�1�����,��4���I�����%�yLa3	��Јe_O�"t1��e�����Q~e(Jf
8gj1�N}������R�t�GD�젉���c<�1�=��Ua�qR���25�W�����l��b�A�GS��w�Ǥi�(-T���Uj2���k���;�;z�X�j��	ӿ��avU�8֬����!������uH5���̐�Ӗr�)T#���d툶g���U�uJ�����C{�D	
�	�y�T�̵�)xu�f�V�oʱw�y�s��}C>��2��w>)䡽t����ȸw��B����Q ��B�Iߛ�`J�H�C��k����o��@�t���=-�uO"c���)�5^Ny[�C��Z}����ʾ`sg�4���PkG��)�_t59��^���36���f�����G�� ��b��B����'n?�8����P���:��>?�>�B%�Gj?�EW�s�KR|����	�xT�bCa6̎��{.�����&�O����|��3��x�6��9���8�)🐖��A	{�T�v��u�U�yB�J3�65j0��(���h5r���������*zͦuֹ����/Ʈ�]�+T_p�Oq�)�����3r8�e6�~��<����F�]�Ql H[��� D���இ����O��������3��v�d����)�KT��<�3�_��ge㰦_/x��P�	��\'	���(��x���G��q?�=8��$b�s�a�Ȇ���9���='�ƻn���@ȳ��	`t�،����J>$x�zB4!�J\K׭V�t���C��j��if��B�)R�q��T������d�稪�T��͛���I:�p���S�-.�=���2��8�N�,7ۼ�%I{��{��՞��93(��4���VE�r�~G ge֐�l_��F =<�I�.\�J�w��7���{�
�h�Ǫ�]��@0Tnj���U����Q����_�T�㊝̥� ���H�/\	DJt}$�2 � h����6a��9ycv#&�ێ;g��!����ʃdn�tiڢ�({�A��Jp�^V�78����g�5�vٍS���]d��k�["~� �G���R��ME�ը����� P��R�.���Qq�.BSlxzޚa��϶| �р�P�Y�
�{���&�#'WE��z"��pl�t���ک������Z��x�Ue����tlm�"dOxi�����R@�T�Q�X)���\V�u.��D�I=	���.�[�1�Ő� �y��		6�>_M]x",�0�����ꈇ��Ɠ�ɇ���*�-"��Ŵ���-M��9#�d�H�>�Д�g	wk�n]�y}��vv.݆�Q��x�hBy��e�\I��w*�h�L�P+�	H̴���l�&_n����_Z$����q����=�Ud��x��%U�1����O�5Q�_��P�XY;�f��L�k��������0]T���!���u'˖a�cBq�qp�ٱ��ڶ�}a�^��s�t�[/�@Q�>����F��umt�Q,)S��#��7��4�]v��'oD%�Ŭ4
�	Ѱ�)=*i���9����K�CꉗJ��/~�	 �����'F��-e
4T ����\"��O�-�"]%9���y���%P�v��f�]���E�r���B�G�}���)c5|edz��+2��Z���>�;������Xq�ϳ����nn� ���yݠ�8��L	�����v�6]�qZz�R:���!��\l�w��v�Z�Uq�����p��t2S�W��|s��BǺ��mJ�t�!��l��oU�I�J��'�Ѩ�w��(N݁��!C�X�Qб).��ρ%��J(����T�����Ut6i���P}��e$:�=�uƔN��_�j�eN���&yX9���w���}�ւ�F(�a���y���k�na�.��H����Tޭ��mp���;���0�^ou���!�N�����Ğ?a�܄���~d	\��倖����DXo�Et��ӅUK�pu0Ҿ^�j�l��-b��X�W����IѬW71hZ��71�V��?�ZPo��,;|�K�x��mJWk��/�b��'��uB��Ց�V&W�P^͜2�=�j>�\^�b���8�`-����^"ͯG����R�&�S��
��g7r$L)3Fr��^�E���bS��j��wvȻ�@���L��`��=��fAm���r��W��"���������_VR�nr�ch�N��}_#^�]A��=���ΛY���iy%9n��,L�V��$nz�OJ^����'��Dh���2h��R�S�J:�������rx ��c+*��� �.�����:o�/
�H]��rz�B�Rk�S��9P_6� ��{s�	�8�����G�����Kcn���aP��#u�G�z��go�ﳷ4i�l�֞,^q���;�b�������`�� ^�Q�
v��ؘ\���u�
���\u<½�钁)���V�<���{�����쪭��P�K- 1-���Q��|���*�"���;�=)�&�A�#��&�)/�..��^'7#���_�W�Њ�M�-��x��yٸ`���%�(H{	��΅Ύ(������A=�r�"�x}eɥ|^;4,��l�;ϲB�Z1��F�{Ӓ'}&Er��Q{��+B�[��xgL�i�[o�qsr���C3�Pǁ���B����;����@��
�cS0��(%U���_I4)`>�Q���<��cC�v�p]F��k��D�j =��h ���CăG0�٬�X�8�3��k2!��f�sʼ,���9���(�LP+�k�v��c���0K�Kt͈U�
�G�� �j~g��hGZZ�h�ry?�$�T'����`:�H ��R@��V�����%��`s@�W�H�:�?�>O?�I*�^uv�Q�;x��]hw��q�l�YzN;��������'�@^|�/��ք1u�*v�c��?+�~���rM]��8-D�{<0u��O悻@2��'�%)tP�ʦrr"5*�@�]CV����|1��`}�^H�È��@��M�=���0b; �,�]�AB!�T�CaJ}�@W��H���vp'aK�>�t=}L�0�pu�a&y�$��W����$�r�D��c�S��P�5B5��Ԕ��S���8�`��'x+j�����"�t�_@�7]9��+̤؈kH^�"�/~�Q#�
f��L˛�Dr�])��!�� �7��~wnn,o�IU��㓫�� q��VE�^F׺�-��M�l�%�l�[����`f�� �^3��@�?L~&�g�o������(����F�U�����VA� %Z��rP�IE$��~�,�D�'�\���4���r׫DR�U�k�������F�˅k��^&��sÑ_��C]gD�f�̫�,��Ik�_�W����U ���䤛����W��K(��O$��@�:�p��fw�@	�E!�N�U�%z�놟�� �C%w��NG�k�ӺL���C,f�q?$�Ц1��}��7"I����X�/��>yIA�Cж�^.���>�%w�L`ꑰR$��:�G7L伄�f����	X�u��LyE�؂��;�y����#���w�6�.�Qϣ�r�p�D���!��\l�vy�J�Z/HD5�F�G%\wb�?u�s �v�!����A-^��G(������D�_��_�`�ґ�Q]0�f8�]����kL�ũs�pG}�+O���������`	�>���e���R��iHn@To�A{yd�����Ƶ�Es�n�J/��ٍ�H����(P�}�*U%�~��Z�,���+���Kw�O��tˆF�\E5��~]�����3�|�i�� �h��(��'.j��A]=���@�į&��gI<V�R�9�*4S�z�jJ���x|);<�`CܶW��~��1�<^w�ZR�� �ǀdm)�W;|Ve�E��f@��%���u �|w���r+����k���!�k ��.we�jiKkޓ9rv'������oq������%O��0��j�C�@$�yN $��;e�赍3�ԋH$b|�߫�0�L���a�vU��o��S��d�/>k����E��6�%V��
Չɳ�Zܓ_�����͕h����Y'�$ؙ�ߝ(Ւ�֔SFr_����;�cJm0���=t5�9$k��_�V��,��͉f�k�`:�dfơ8�kL���VՐO��P�>5��M�f������]
K,3�:�b���Α�m��YX�}���d�+�T�I���1�G⨷�拑4�J�^yK�p�%�<>[z7}���S�9	���yͮ�z2r��:D*����o�lXi��ۣFdɠM^-{���̧�xw��e�%����L�0��@l��r���ȴCm�1�!��a���]9N����z��t٭e�7�b���l:�G����Mw��β�H�Ҳ��,���ۂ�t����e��'jL�Bp�E2}Vm��I*M�#��y��>�z��J\�>ơF�w�_�U�=�M^k��F�m�o�����6n�|��ˬQLI��B;C㌕�s�ߴ	¨�W����[�=�Nsg���8���B�D���h�4*c�a,���c6���b5���Rd�];u��<F�m��͐�I>��,U�[�XA�Ld�^�v��O�&*7l�I_b�� �ԍ�"�k��W(A�,�t$�����X�S�2��X��������L��w�x�� A���l��u嵁�+pd�Z�c)C�,A`g�T#�{�Z�k8���w�>�x�ٖ>�(�~���1���96���OJ�ܟ��M$�Ņ}P.�_�����x%?��1� ���2R�v�B6���+�+S_�'�����,�X�B����f��[��B����ތ)�����:����1*mP���{��D��)�2i��,V�v]zÅx��W�;8��Z3��T�-P�'�ۇ��`��@}�b�@d��p>�֭X��d�g��d*f�,HI���!$��"����S_&d8�e�ڧYU�wܹ� t��ɨ��ـ�k�A�|�k�6�2����r���b��G�"�c� ��(�@�#}��>��A�P3��tkV	F_.)�oo'ʚ؀z�X����
��~�?:�[�L���Tq���_�F������K���͆8�53K#M�GС�	���Zj�u ��o��H���/B{�#ip
����uL�\�m�1�
�{	�
E�}��~�>M��{��a���s ��{�_u2g����y�WT��F�D���w�΅�KQ|���	��:u������&N� ���>��u�j�4���J���>&��'�`%�2SL��+���������0��z�IM����]5�3����#�x������3ɘ+��Ϗn~�_����e�%WЏZ0�*EmucJgp�1����&XY-��fu䚐��lc`�����G�&g4&�P�_nx�y�u��)���е�'���Z�̺��v>]Y���¡�E��e�
��$�O�q�ĦK�p
c1w6hi!В�6L�a�!�paԅ���cIH�"���E�Ŏ���WUD�BXQ7T �nR����h��0Q�k�����ĵ	�+5��	H�-�|$"m ~DƉ�3�>v﯇���2w��5�<V��|�K0��a�8-4۾ V���������x4�II��!���y�.�cr��1G�|�d��C��q�B��k?�!����{'���{����1�$ ;�W��推Fi=W�*�+AE#�KA��	���]&��6���&$_~_wN��90bf��k-F4 L���^cG�*�Q��e\o��h���n�	�F��A����d1���K�In�h���K<�~��Ƣ��"\Kb���� ���~ڋ�3�53�j��67��~�� ���͇����idd}fS
����%9�o�����=�|�h:��j�r5�[m�tF�KHh��9Ŧu.w������u���������P��FOw����z:���T���Mm8%;�;%6��O	�h��˧�����{6SXL�gq5ctA����� c�%���H
HIY2/�|�ᗴ(��j�Ϡ��>�Q���}FKl��1�~i�XΕP�ԯ��x��WlH�@��q��w�w@��(~�Ui��{7J��0����q_TIÆN"���F�I��I�B��5����o+�J�2���Ȝ�h [0���*�)7#��l���b�ɕy�XJ5��Z�b�iq9*��������u���5�,��Z=+q4���r5�$�ɇ��6�;������Щ��U<����u�X��h �A)>G�e�MV���<J�q�P�N�������7��@`(�x��+���sv[�_N��?�f�e��� �bX;�Ɣ���I�����2����E"L�|Vtyvf(������~4��̻�yg���v�X-�[�Z��/dܡ��%���X�{���`U�G���'�*���^���s�V�2@�D��YG×	>oi�,EG�ŔdZ��K��
���px!���y�	��>%g�]C���C/�ħ�m磏�݃D(����໨���8ӿ�`B�F�G�^���O~J�
��q��/v������J=�Ǜ��n�hoQx�m��s+{,����L����� ���p���F�+����S?��TU������?�V�x��~�D*Ae���ՙ9��ޫ�p�L�3����vׄ����-�&������\��9��j|��B����^ ��I��WR/�t��=�ʮ��6"=���Ǻ��]	k�vO��b�!O����f��!�
���~�~d�L��9Nn|�1��M	��Jue.����j�M /j�<�Z�E !z�Ū�?eI������P�nŽ�.�lߔ����l�,���"�-�v��z�6�A����C�u�0�upT;S��Ӑ�B,�����)��n��ml�c��q4�@�k���m!���7���Z#qy� 竈���~��kF�,���\|&zt��8Z���� ��M&�d���ƒ��4Ž����w`RC'	t��Xk��g+D�P�����8 mR|N.�(W�	F֛�cᶂ(���t�S!E��o.�"͗`�mk�S�}�KW���M��+�2�ʶj7�zskO�=���`� LV���.$cFO����%�ݱ�4�9�ՙ�5{�W�������v�R!�ܩ�Ӷ׸._�He/`��2t��h�cB?G�t�� �Т�����|�YN�/A#r�V�R!Uu&9f��.�N�dUY�����	Aa6<�Ic���])�ߒvfJ����/~r���Ke���mJ���P���!c��v�ZO��˳