��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�oA��J����� �)���SyLw&�JD_�,{��X��%2����]��FJ�
�Pw:�>��C����S����������j��FE��xod�d�/-�a=ū��y�,�
K�[:�iu���0m��`?`��a
Z���*�WF*~2�$��{�+R��Aꇊ!L�����+U=X�C\�s�.�e����5u�e����}(Օ< ֧;g�3��a�������$���i*���ɪ"�qRqP�ߚ���ߩ�����ZdL���ˌo������n�ڡ��O�>��~À[M��:�i�Zu�	�����А��b�A> �����~a�3�.൥�׏���=#B}�؄��y�vC��}e>犂G���ث�����۱�8��ʙ �+e�-@f�W!8��( ��d�0���ea�V�km�θ$���F��Q�Z��B���;��^?J�IKy�K�M:���Dod�eX֛���a܅D�`�p~�u#:m.憮���i�2����-n��=��"m��WG��Q��~=�jT_=p��g� q�)S�_$ �6ݥ��b�&f� H�ڷO_�}O�K����l�~�rBL^�?Y�;�@^T���,�L�s�ʰ��w1
�X:3�E��>���n��J���r�d��s`xdRk����2�\��y�^���;EA�M8iAAJ���M�{���^&��Ə��ZH����԰L���!�d�_Y�V�&-8��qKЛ�xB�e<�I�9W�k!ɘ�֡�cXmݮ�s�	MW�:�K:�o�F{�(�X�Sh4��KZ�wOJX~��y ���}9����oaH7vQM�QG�K�����ٺ#�<�W��L�1 ~c,����چ��-��ɔ��Nc���L�g.�'�}=�l�$"�"e��s�1�(�|z�� �V�y�({�s�i]��)o��+[�cP�ք�n���lB�]q̞tQ�����#3���Ʊ~&��ߴ�0���Q��iɄ#�Z]�4�:��7g��7��5��u+�5�Á��З�b2��o8��S�2-���ʇ8)���Rs��L�j ��=�ە�����a��t񡊧m�T��G�O����x�2�)_E!�D�avP�=�t/ �d\��F�Ju�Z,a�QF����G�`�%��l��!+)˄;���d��A�*�nw�\*��n��m�@o:R-�� S����g��j�ٓ�Kq��8�}�*�ʟ{6�>B��Y��a5�;}>т�� �I6q�Ch��2�����HL�A���X.��MOI����̏��êC`�z��� A�>Oa�+��;�p�H���M[,W���v�#,�J�w=F�+b�!�(޺}�C/_�S.d�_3*����ף�S����NJ�Fu��,U��.���F�]$K|���j��r�#;��o@f���Xl6Ϊ�&zb��oy*�CrC���&v�R��hW1����J�{�R�x�a�Cr�~\X�_I]���Fw��1b'E�Tu�F�~Se����L�>�m���W@� �V���6�Y%����a�(#�+�<-NC�4�{�z���d��$|�D_��$�w"&i��r0��Sϊ�<E��Ƅ4�׌���0p)�y����Y��,�KB��%�CAÎ'p��g"�r-�/n�[������gd1��Y�?��{�`��tM���!��A=��uԳ�,_++�[�������4tzY�]�=�_�g
����4��47��|&��T�����|�K�n�a[�fV1�{!�C��6SɅz�1��b��t���OS@�� ���IA�_eq��5C3��z�����9�f!pLҐ�kj/f�M3~�ޱ�݋U��K�Ǡ)n�]��b�9�\^��(C�1G�7n��	L�s8�@�=�I�����w6C�"|{��7���T󄂝��2�Jɼf{�}�%*�D�{���g��a��Y)�]k��]Ri[L��O�c���JF^�f��tr4S�m�R7���ũ*fi��*?8~�x�zQ�Li�.dz?�8ʟ�9�
��ӤvN��P ����Ѻ����,Ǔ>�����0����U�Cж����F�E:�h��V�	E����N��iW_�G��j�饯��n77� U��n�-��8�;�h~~
<���d���}xn�Wγ���*��"�d~=�NZ3�w�ցT�����Ee����z�[Q��2�\Yojg!Ӻg����l�X�������@m�N�-�y����lD��d�����q������v�А8a�eig�^��X��Kak�����m:չw�!��ev�%S���s3���.�!\C��;u�I0��~(�$eTu���sc/�t�l}�M�Ky��rq9	��fG���PL��	����]�o�+4��,>��vv�nN�]��xz
�$�oL{�P&_�2{@�"�l�xR^��l�^Ɵ�˃C<�㖦�%Y��5�}�Ë���HV�Z<J��G��8��,D�=d�g��r;��������O?�	5Y�,lr��:i�}4��(~���H�T���q����W�y@�= _�cp���>d���-��`�©u�ς��Y"Z���+]���  M�y\�ļ�FR���q�M��q��տ�9���E��q��I���pqDN��FPw��#�Jv�[$�"��i��nf3�{��S��mHϳ/+v�ܢ��B��˗�%�2�FQ�~K�N�5C��U�CRy<�Ƒ���7��`A� �����	�F��v%W ��% �X�����n}���w�O����?�����I;��¤�51��Ɏ�5���"��2�F��U�d���+�
d�z�TGxҮJ��&m-��Z�.���S�I�@A�A�)�4���,�v�42��] ^�]Y�톬A�N'���.�t�9�m�?��q�LE�)4�z�;�ȭ�P�:BM�����l���6�����!�)�o�?ruF��mU��ɰ%��g�S��f�� �-�\����̈́H�մ���DJ�w�㑘.��l�4�<~���Q�+$0X�(�H�
��e�ci(��ܵ�Ϡ���6.3�[���+t�B�$,�p+格rc'���Z�z�i�le�`��쵰Im�ࣕ��>2*���*e7�5cd�㿔��"3�?6S�0� Aa�<��~T]T�jV��i�הAׁ���&BЯ��%=�����,�3�K?�E��z�Q�WJPm��\�^��X�Q����u"t��!����T�}�e�4�8�A���I@���ňJXz�;?K�jp��A����]��gQPVd���.h��eE=` �u��Q���*�������/3�u4��g�؏���������}��r|��'<d��۟��p�0p���9��%���M�J8��l���m���g�m{oW�c�`� �[� �E��0{�8<��~�����&YIw&	�Wf��-��E�Dvj��Z�ne�l���V�0&�� �Q,������tZV,*c����܅�#*$��b�SF��2;�U�l���2Q��-ҟ�D��S���Ɇg�T�S�G�r�B���v��}ҩޟ�ʧ	�`A;-4�c�Ű����լ����}�i��A�uڰ>�aRmO�N(�ґv��`n���-`԰�2o[�0P��"���/N6�;!b��ҁ��4�#YV煚2��;��~ᐭ�>�u�b;U� ��d�_��j*���E�W36{���Tɞ?12�fs'} �7[R�l�'z����巴��6�泯*�~��t���Dr3���=����KiӍn/n?糑n�	�4��J�O*)F���sd�B�hI_��v��s�+�ٜ��隘��k�*�v���i��0u��C�Q����͍�U�C�rC�A���/��:ͱ�`/MN ����
ɚ�7����T;�����p��!&����󲥗�)X�ީj7P��Q쪁�$'mc1�
�����K(�{^�D6z.�ck��t�T��3��cB1�NAN��e���"K��@�I�R������x�D��Z��v�BX�Z�T���9��TN.k�Y��ɡ��*�����	6ۀ\��@{�7ɍ�H����u	��ޭx���j�鱱�E�/�A2�Bp�6|�E�5!1�o�\�s��o��rf۠jdż6�$p�G�_!ճ+��� ®�.S�j�՞ï��b�D��d��m�6���m�b]�3b���䵥����/'P�v���l��κ�S8E%;[��S[v�]f&�pב�������6���5%K�7�\G����N"͔���+m���1�kQ�Omw�R���H��w�}]��1o�o�NF~�)y�F'�;���t������	mJ��A
np/a �{��P����!C�/#���O-�7T��T�lJs�Qw�w�:y�
�.Z ���vѺ�t��É��8�q��Iiv&�t-&7[ f��1�ց4�2ڦt6u��������������&��2\+M-�������E���sA�i�3�9���B�L�+/9�����cq�`�/�6v�9z'>��� �Y`UQ"��P��S��p�'za�.T5��� �)�x%��`5���).��iD*��r�ð�ڔ�<���a��Y��~*��%뺩�w�I���&��*6_j�V������7�i���{�~����f�L��&��6��y�=#w3�G��|���B��$�`o��������\b*�����`��T��꾤����۽�x��n�d\��x���!"br�VS�7�N���-x�)�\`[��@`�[U��vD��2@n��
�WC@���l�Ϸ�@��X�����XE�1�k�I;��+u}}ׂ ��NJ��+��l��5�7o��H|w�w�ѧ�E���碁�r�t�8U�{௲��A���@]w(c�(.�f�;vp����yڣ��H�~x��"�x���r�"@�L�%	&���y Ϙ� �vI�e�>0]N��
��^4C��H�Ձ�j�^&��'�,w���Ʋ��l+����\�/W2�?:L�	j�y%1<�}��x�f'6K�\hoRx�8;��p��[u�j"A5L[�����3"��	D,ݗ�	@N|��\�䬜�K{��C�y��Kv"*�"]EdJ��P禾� N(4zo��l����� �Ez�	|�$|��<��t��|{]���F�/���%��Ł|�x�x�N@�,Zp�)�bl�XO)S�Î����i���F���AJ=��G�~�4	����ċ,�\ �,[	��|�5'���%ܤ��"ͨ'�"�s�(��� 
�s�_H�~16����Q=��"�o��4`�S��rMX0�9���⚶�S�t~8��{���a�^���U�<\�����
@A�N&���!E`=���z��@ l�hu�+1���%2�K=�"��$G�p�
�D?�_E@ǣ����� {&�H[5���5�r%�C���;]���Xs����&\�;�;^�;a9�p�,��������U�������`���˨`:�=6E�Ç�tO��h/�F@�9�r�>�V�A_Ű4s�5��e�;^���[T�$쨨���^3���K����Q��*�hG�4n�BߒJ΁��R�OZ&���ME�ƌ�$����xB��Ƈ��,#GwR�±�7쥻�\/Y� 5�'��w`��>Q�N�Ns�M��/�\8q�6i�yݴA��ϥ�uui��I�Œ�(��a٘Mo������K�tD~ݓ���IZ�Cߦ�w���rW[N.k�������B��]�:�\��+��Jl�[�"J��0K;mI�5��t��Z��O$���N����q�c�d� �0?��R�;o��Y����m �#��/��5���BT��d,tؿN�ʂd��y�M��gE(�!����C���2�*�_g69��j�ے\e��Ob��νD��A�������V���jR*�i�M�Y���;�̋�
1���|T�+0
�*0�-q[������^}���Z�M���(?��?��w����x-���c�f�b"�e ��F|I;��s������OI)9K��]�d8^+�ٌ�������:����~�>�5�^���x�3�*8ē�F�~�N��lV��8X?���ᣂ�5P�FA��"�r���|G��j�Wm+����N��v26�ECD��׈�43�&��He�8me��viA���)�V�3�N[��!L�ɓ�?Y�o4��eAO����W�0d%+1����~���嫲nJ�=��QtO��B5�I��)��c�������}��y8ώ!�H�q6��	S�g�6�<���4J~����$V)����(0��T�3 !5KC�/����$���n�n#y�Ϫ3��
�� %c5�m:�Xc"�0�@E�({T�d/]���6��=�R�c�Ϳ�M'�yx-�d����%K<�f���V�����Rr�m�o��
���e���
�q�Uve�Q[�9
�o�Y_�x:B�CU����[�t7S�`���rz��FcA�Υq� #������21��e �w�D�},� \\r��r<P���Bc`��ִx�8C�M|��]*�	���=�^�W.����i�Ĭ+|��ֿ�ɖ�%6Aۈ"Pq���q���}J��ٕ/��s\z�Z8�IL���Q�uě�7�������2bM��~R3n(q�gu8w>V(�؆}P��M��4��\�=O��$Icx= �>W��&��@���S{��ꉾiLMPĹv���Ov��(��$q���]C�:�s�0۶�~��1�ȆY�ݣ H��׮�v}1��S�ym�ǿK0�~�o#
�T�����R�߅C�L����Y���=�	��D��y���@T��-������7)�dϷJ9�!WJaR�G�98,Cz=�(��sU"bW!ii������,��G4���SW�f�K&�~U +5:4U�M�E�}�6�l��eXYŘ+����"��3bچ�%{����	��En�r��n@S�BS׾�}��QP��t_/�Ȓ����.+8+o���w�L�h�V�|����10ؚ��G�8-AxA/�+F,����q�6�nv-	^E����֓���[�����-1I�Zl|��|���9���h׺ەi�Ժ6zY���d�iy���-�cw	ֿ7����;{k�Pw�����&�=x������{�K�E�U���#"�+Ȫ�= �@�:R���ԡ�j#W
��1!��K��9��^���'�Yq(�ZU��|+5����3��E������_��<t��g�3�e9�N���0�i�4b㌿�ޕH[�v�
u��?}QZ'��<}��R����im�gs�T�2�Y���\R|S��ÙH^o�@������>b��I�%[yؗM��}���F�Low+a��y��-���TTi��A�DE�VՋb��@�/�۱��/^nŇ��EJd�Ùf�š��uq�當�Q)`|��j���5�4���nx' _�Qϋ�4]�4Ǩ� (��[�,a���'���bQ{ s@,�ѝ�(���Ÿ�$�3&G��c̓�P�=��͔��)�n9��[�������P#%�H�{�GoXb�?jݗ5M��_��v��膖�S�Ū��P|Y�$��5*� <��e�Il6S(-�Թ�^��ah-���e3etUej��v:[��!�*2���fIt6�eMf�e֏TFh��K��vmc
�g��Wݠ1u�Ԑg��6�-�-�
R-T a���Kv��w���Δ|�/�(Ǩ'|P�[� �	�H��sZ
�a����c�Z��.瞒��w|Gw��$t:Bҗ�����{f(��f�Ԁ~�¡�!��Q�z'�Q`-���CÍ��LK���۸mdQSj����Kr���BU_���إ���A �mp�@޳̈��x>:'����eq���&턻26	�2��Ͻ�2Bp���He��ݻ��:}P_J�S�w����6�P����s���x�@�8�m�@ũu�S�q��.C6f-���D��N���gݠУ�Ok�a�N��GCP=���N�ףP,!��d*���7Ϣ�&eW�����9RW"~&19-���� N�Z�����7wo��BM'E�����{�o>N�"F����Ħ�:�`����(R5���'��W���Z�z�c�;���G�ap�|)��m��U�#��L˩qȶ���@},֙EP3[S/��&T)��销R6^���bY�+%����k�E���u"�c����P�M('ԯ
޸��,���]����BHo��@twI�!�N;ۦ�h��cÐ[y�!�<�2[t���J�W��/)�h �f	To�.l���h3�dk���q��-�(1�U'�J�/�&Ct7�ez`������{*}�R]ءLí>�~K�~ ?����0��Z�t�0�vE� ����~I�WzD���X�w��T�		o�4�ax8VO�ڸp��Ml�r�=J0k�R�	?�> �qk픹U�#0��ky}�<>M/݌l��$D@�Kp�G�8���E&�r��	�<�j!��Kah��{]_��"�ʹ�MF��?��u�J6�&ت+�U5k1�N�������Q(|،h����nJGp<J?pZG��k�@=0i�ǃ|�4F���B
������}zQ��o�Q����LdP��t˧P�Xs�a�J?)G��J�)7�z�9޲���{GeQ�{Qm�����@���-m�V���sY��ڒ��yC��|�f|JjQo��5�z�
�ݷ��HM��-O���D�h���ׯX���cl��Z�s�O t
�A;�p�L \鿴��_im-�(��VoW�����IR�/�]	�-�B�є>��h��xВ����Z�p�jEL��&w$�qq�>�([�ҍqx���SGȟ,��5DRΡ|��AIU���4p�;�=����� *�8�^���[��$��rd���*��q?�.O*��^�G�@�ߟ�®�C��(��.Qʚ���mok�)Q�(ѯ�d�d�/�<H���x*Y�S-�=���𫖡���#�B�8�x�_c��PC��|�V���R�4� �������79����3�-��l>��u�T���a��ڍ���$ߌe�ʍ�7��1L&	n�ݠ���ё��C��[�,x[ �x=qj��ςʗ�#�M���B{!���gT��t7^�Sy��y�6���j���ɣm����?������+��+P�1��F Znb��"�jC[�����
���eM��@��eQs	�㮏J��טPW�6Z@����������Rti�n�]N�7 �-�ʬ!� ����xy�J�����/������ƥ/3��n%4m�Kgvi/�`���G7����V|����j^��;��VA�S�T��8���r�i1���e@TUN+Q����W��� �hY틶D��CD�����TH���t�E#
��f|z�tp����(��+v%s��$�m�򬏆k���<�!y/�b� �h�${*�n�H�`U�\���qW'��J��S�(�X\�����!Ob�����2�4���I��̃�\��<�����,��c����d
��`�����Ÿn��4ʀި��5X ��v�{}�A���41n�|[�+�d��h�%� v�$B��V���g;3nr��aoo^������)����_5��I\�z9	ˋ8�K�cTd3�N]�h�.O��>��25f��2���1�5�2�|Ū�'��֛_�����-�ڙ��`0!-Cn�>�c����f.��N��`f�IT+��|�?�.�̕�7x�|��=6DW�X��7h3�_y�_��K���=�t5ɽ����
;qt��7,UD+�U���Tf�r�����C�q�n�h�BJ�$�M�� ��(����J��K˺�V��Oh�/����'J������h���_+�_b�V/$����������;���,��J��=��9_��
f�$�1+B ��'�-w����X,�B������A��(��/	z�J��)T��p�����A��%���O�:�m���Q��繲1Uɼ[-�k�E���M$�91�9�4���ǉ��������(�� ���Vo��t�V;�	e�P���[�˂v�����������
����, �^g�/$��Q������O���A��<��k����l�B�E���6!�����ؾ�	 ��%���)���.�j��X��X���Ff]a[�p�363��'tۊ>�	�C)w��:�+g��K�+�R��q�鎼T"O(D"|��ܛ�d�l�Fq?t�bL��pڄZ�Ӽ[� 
��#CtZX����zD�N�YZ�mast�S�Q%�����'�-�Z&gl���S�Z�n�X�3���8n��&),��0�|�g�')�KT��v0Pd4�	/8BNAT�~g�� $�zq����ú� -��n^��{�1Mt�'I��p�����G��<�Q{21��G�#}��m�QI���`��{���X��*��(�B�O���3QL^��R��L���u��-���%��J�-o*I'��x ?��o����� ��wS��N�0"��~6�(��6}4N�+5$���j�nH�݅�nP��O*�X�5��xD���o;#t��pd94X�Z��g���/Ie9mQ� :�;P�K�y�.��:�{Lm�wR;���l���.�V�0΃���l��e[�<�9�	M?�C�d^�/?}�;����b!���@����f;�Q%vЩP ͘�c��3�ⶉ�=T�,�eM.�P'hd �Suyw��H]#��@�R:*$��DQ����q�r�6�ԽbuS��;����k�c6�$'ō�XtcR'>�7{
\�
�"M|����$�z�p���u�rRܡS�2vJ���K�����P�B�G�W�|�7���v䀐 �*�����3`��k�8��>���%f���8�L�8(PU�[]��O�M]�*VKc�y��u�F#x�������Nz�	4���ڑ����Ipsv%�h�&�*��"�L>GAv���@@��P�xN�.�<&;��S�u^y6whh�nw����5�_΂q-[��e������[h껲;�w� ��/O8��m�qY��¸�x�KȄ_@ro���R�MX�A M��wť�O���q,x��BG9��P�糷ȗia~��j�`+N]+�悹��~���TF7��;��f]?�=�!�������$��HZŸ�0%<���H����#m��@Z���E�
Sa�]�<7&���(�A������F_l������U�Hb�E#&��qX���ő?u�����a���u(<��y�F���<dCB�s�gu�S�,��F�C!
�[�Ա�<}I�x>��(r�:Ud��*�j81����(��	{����\��h��QLXwJ���)��]�������\���d�j��,r�����w���+G�(i��Y�U�{�/��m\�C�$�Q��}��(������-��S��F��ڡ� N
7��b��Ϻ��ג�]hi
h<��P3W�/@�e|_��t?����{TO.� Y6m@����o��Ms1���`@��]r��h�0ua�� �p��.�Fe<�OS�Hi��3�Xr(���A×�PYe��tU{9r�RBua�m,(�4��$OV]W�ٽ�%�S�fs�U�U���J��r���۠ �7��W5�t7˴d���r;��� �q�L��<ۀ���9Xۄ���K�Â�b"u�!�%F5�/�2�4�Aj��G�����X8%\N˶����Kc�Q}l�{���7��s]%?��u��3c���}$�x�N�Q����ɸE�(��7 K^3X�up�"_)]���G�����mu`���T���C���r�O40:�����x��5&:ٔ���ۑ�'�E��-A�'3���E�9&�×Ե�Iܹ`��M��x����<hf�z�Lr^�Z�\��4`����c0�o���7Χ�{�A(�΄[pč`x�YV)8���Y�/��G/Mr�os��}��fFqs	Ü��U��0����\��R��LE��b:f�TK:���⩤k�!KfNF��
q 5��^��ϼ	�=��;ř̴\:���O�<�����+l�0�d��:0:�f�~~�cS��+�T�>������=��.�r���<����	��d���]���%p��]%9��֣�x�s��^:��,8�h��,��Z�vC�\�<j�7Ņ}a�!�}����MW4�m�~��K��+=Lڀ{���ӯj�֞��K�r��j�z�D�'���N�F̀�l�.U���ò��R�=����m������M1��V��4٩d����J1��s.ܢv�#�n�p��	G{����-��[��&�-�#�"#���@�����X!��x�נx1����"�0R�������"sp�Q�g�(���t�Q�JP�6#
Bҕ��Z���ӳ�a�~2�,�e�)��M��)�����0/��m!�R/�.��򑰞°*h���@rv���qX�$[ @��߀��t.&y���q�
�v���wǐ_揥�K���Y�>"ݴ��MX�^o{�/�Ï>sw���egR�(��?&.V�[Py���t9~��3�~=2I?��b��,����2ߨZJؾj]Mk� A�duϼ���DS&әG��34�A#�X��7I����$<ͦ���d��T2
��Q��im��tp���E�K٢�q���W�>�|ǭJ��~��>uo^٦<y�.C�yC�j�N��S����,�/�@=4|J�6�� ��Ȓ4zY+j����N+F�ʗ0lHj���J��ks�˒�O�a��M�hLXs2_J��i4��	���/}���]��	h�wI��9^�@&�o�QO�\P�1��=88��z q2 �YD�=��ܛ�Ħ_�����e$v��}M��~�$L��l�K���`4� ��&�`��`��l���]����r��ʒ�-�<g_�d��AD�,�xi�8�q�-nOQ�_g�iKe�O�Ț_�(�6�X��9�$��H���,��'^9�'VL���k2��V�b��N�Iv#P�(�[t _Zg���v�	"��7�C7�a�(�+���J���ˈ\F�=$|�1�[���Ν�����5�K��ݎ�,�1c�g��{:�����{�4.#B��u颊���{PV.y�Ռ���`�m��%�i��Y`��'"18�>�s��G3����8����ZM�
>R��y��%Ռ�����5�k�-Qr�\w���
�gI�47��1�x����8'�ȣOn}��uL:۩3�����yq�μ��|р�-��J"�f '`��&�QE=Ž#l������+� �4�ن����N�h�`���I�D��D�G�#9`��㺙9��Z�+��ʙ�q�)d�~~2�����Q�Ü��4y�_����;.�f.U��'���*\�
�!J��t	JE������e��F�wY�{��O`8v<-%FAа*,R�}�۔oV�(�%7хHǮ\�[$��ͤ�E�&�,�B�\����
d=�m�̼��24����-�|ݱ]Ves.�ug�����x�	c����V+vO�J��.g�Wk����a2`�V���4'#լA��S�����4#S:�'8����'@3/��㠆� �� ������^�8b���e�&m��� Ό�}����`.�߼�`��+��OS�W�]����0_��)�KZ
i�P���5I/�C7l=a�u��z	�7�Y84R	.)m�(cc�C�}n�m!��4�H�h�_^��*��9�K�3���+7�Ə+�t��9j�,�g�ٛ>1"쭂;J:����7����o�`��J����B�1S��t)#Nç��zfY����=�G��-B�?Z���y6On�y��������nimu���fl���U��������=��h�JU:r��{���.z���M?��b��N�f�1��75gT���Fg ��͝"ԥ�.Q���N�w�3���'�N^���t>`��h�Z��;6��k���K}$1�I:�������)O�J��������Ap��,��HH�4h�΍�����*'�Q��'�(`1��c��)����{��͒=%s���q�Z�9��?&��3`�]¢�%|:�"���Wt�ϲ�|��{V���믷M�EJ��L�S�[�Z��+F�0���6����<Ma��l�����?��X[����r�1V���a4�>H.eN����H��ZdnH���ͻD<x5i��U=(����r	��Yy��g������xl���P\P`SDY�S�T�0(��-3M���yS/�L��qr��T���_�_ �a8�`{�GD/}S�n��A����T쬁+���G� �"�qB��eU[��;U%JYі�Sa�	O@a�T�&_])cJ���껄փ��nX5j�@���o�~�G@A�$�ȚRYݧh[[MC>�tpx�������w�Qp�o��Ti���ןK��L����Ň�<�%`o�5T�Q�y��Wa��3.��K�r������3
bz�¾�A}(!�'�R4���.'����v���SZEMB�
|7Ot�B�b#C'&M�NZF�}zL�\��X���^��on�*�=�?�`�7��{A?�U"��rE<EG�q�~5����?�lX���8�|U�L�L�N�gQ���O�߶ o�Z/����.i��(�ODѲ�+u��9E��w8"b�n)�Sp�Nwjm�\Ƈ���&j�o�Hk�-
i�5X�V#EC�������v����H2�1ԕ+�{N4%[RE޲B�	�D 7�+�)]�=?A��mP>����߉�tz�oe(���gP��l�ۓ�r.Ax��~�Ⱥ7B�Z�p<����|���Ɯ�h8�pAw6���5�fw,e�s���\� �=�$�>W�R��Kf���~���q�1@+E4٫�k�nȋ紖��b��ߎM�	<�G��QDt)O��B��d��v�$B�o^��&A��cw �X�����ژy"�(w��V4[�o\�`(bD�Ьa)��y�ٶc��.~s���.�!#r}�xPʆ�!�9^��6V�[$n�x��<��\�}�m�d!���@�*���}�\s=ɏ���E�$ÁI���
vUn׭P��!�Y��G����Rݹ x~W��MM��X@��x/��".�2S�^���H[�̡N���9\�t�s��fN��o�r�V�yY��z�n�Th�8ףZ�w����sG*9����F�?�����A��d�Ч��sUR��� �'��1pE��[`3�R�00�]	F�݅5��h�Rd�H_�'6WO2�S�@��?5w�b��P��V#�OGH���a����˜��>��QP��^��i��٬X�5���@�h�=q:�z�1�C���3s�?r���$3�!�yηo�A,�tQ�Cl��@%`]�S�:�qE�5�Я9yD/5�n8���F�T�T���v�w��_%�x|���5�<�rν�&{��B��~t�hd�@�%�j۪��$/؎5KF�j�}�S�[8���|������;T�/�1_K`�H�фK��w���D��%�hyz��M��� ��
�'�5���\�N�>�}���	�v�b��w/���rK)i�4F��؝o�֩?�%����Ԩ��9/� !<�%8�}hkw�I��O11��-��S����DL�@��N�ѫ��x2z ��ỷfܿ�6�iώ?� �n��n�p�K&s���khh�+��{�����	^n��q��d�s<U�DCޒ�q���Ů�Dol�@�I����M���2��s���(�v(r�xRӉ;9������t�u�p���E[M���2)��||��lY���c�v�����`�/�T��Si��¡xʴ����ء���!7�8j�B�D��ܑ{uiA�����&���ۘ��3�F�T����b��>V1I�b�x��U��t&�`�~fm������ʖM(�_������]bz��u ���4������@~|G;W=^j�Y!\�=��o�������|��1��3_��S�Ơc�����3�+��!����Խ&�|h���j�s�ͭ=5��b!����mzD��'��3���li�.�B����*a8������aIӥ�7����(��\'C:����+�S���)�8��ө^u���$� b�(K��iQ#���'�u�&,u����'Ɨ��,˕/�������AW��3��;n"F	W�c/E��{B-��OA�ޢ,���yv�T��n*;/m���ң�o�̓-���&�M-�[ߖ��b����*�%ӖŞ]S*���Y;�=B�c�����%�t]�N�e\~;0�e�ݖ�41Ԗ��Y���p��� � ���\!p�!���M�-�V�x62�>��w�F�@�����ʩ���=����fX�M����ƫ���w����sV_��yO����K�����x׾\7���éț��:�I��%��x��Qg ;�{���1�|뉉,\ֺ*p������O���W����w��pq�a^�qfnU�"@��P������D��Fe`�[�R�xP~_�x��(C1�8Nh��_�s�Y�Zu: \4��c��Ɉ�|�Zf`7O�_�= �̃�jt� "ێ��?fgw�:���H����Ԧ��n��e偅o��8g�rdk[Xq}z�X.qm�X���A�t��FR������+�	�S�Q��=b#��׾��Bo�\LA�T������L�$v}�M�t�ۤ����KB%:��H{]�|��3�ݍ�MPTft3?}��t���4�YZg�2��Oƾ�5�l��E��q{u�����i�g@��FxG<�������ꧥ�ݮ�କ} �YiRk�hb!��J#���`����Rl�����Ʋn�8�d��,�:qf8ß�9}���.����K�^G���8��w����L�{�>��8����4�R�ǣ�HF��]��U�>���/���/��[́]z���e�]>x51�I�������W��e��M��VUH�g:#JY��+T=���N,�aUp�`��������� ��;�6R�fc����ᱟcf�M�ѱ^�Z(Kyא�b����s(>�m/�tI���в|O��J�����>b		tx�J*v�#0_�@>}Cz��S�ꗕ�ְ}�����@�O)�Q�_���ᙉ/5�F6GC�<�׾�J!���������iyz5�������D(n=����j�Զw: �B.�uT�K��AbG�(6��e�a`��wDI�x�N�b.��9�H����
��K��t�5�rwt��BP���@B� ���
!+G��wj�(F>R�RS� �jPѝc_w���VZ&	7����(�]�~V;�Ӌ^���5����5��'��H���;Т�Ü��P�"�\��^��.Q*aA�v�uoN<��#F��}b��j�JFM�Bd�m�G�=�Q�Ej�*��ͱ��^u���3 L��G�'}S6-*��Y?�)��cژ����X�R�R�_�^8����7l�c%��G���t�f�1��W ��U�e�ŵ�L:�������7�����E��
lpB�7�?��<IҤ7����4��i�6����As}H�i��b	2Oi���.D�m`L��0�i��8�D'���v�����O���������y3���¡��I��ϡ�(���(�������uyL��j�~�ik��� V�In C:ͼ������]e�����p	�m�`e5�W���>ZX��C>��m,\���� X�@�%�;�f[�+�B�܄�mи״Qc���܂|P����1r���6�tW j���PT.������k���1�o�rZ��/q�lm��!>j��aKy|���O`ųQ�\�&�=�w�گ��bw"�|da��|�j(d�X�;l�Pb��ދ�Ť����:����䋃%UӇ���W��H*P���[٘��j�I�p����_n��B���|���9������MD~��ac��#����w�ξ���p��^Y޶j4���~c]�Ĳ�Y���#�E���ى��`�o �I����k��>����#��7�Iz�ԁ '�u�q�B��9Ρ�.� ϥQ!h'���ܡ�+�9�2��3�rG�̕%�ܵ�o���BF���� ���� 풸z,�����S��3�V��/gE;�E [�OjƧE}�v\�{�a�O��d��A[D��[�������/7�g��^ce�ߧ��k�-�M��Eqa���'}�� 9�y�B(��~p�3Y�h��Z���� ��Y��<� �/+F�9��$A�l^�8��&����`��i�C�:�[{��(T��J�yu�m�Ly�r�Ǹ\��D|p�E$ɕ������i�~�,�	\Uz��i��,ֽV؀[�:a�����l�^L[�|R�.@���d�T����V�����EƗfV"n�h�E7A����Qc覶0EϢ��K�����o���F0�p�p/���f�	 ���66�v,�F�p|���BW�"��e�(�!�b=%��P��o���	=�9]q9���uR�A�W~֓U%T2�x�_i��xO�yf1B�8�,iש��h��McR0;�d߉�="����&�F^Q���i�W�E��j�K�����Sgφ�s٣X�X����J'q5P�B��@��-���j߅�KW !ƌ)�ԫ���V�wWm����X�'_����O*!?a��K���Ē�
�zb�DFX���R\`��1-uCL�¬'� P}�2�	Qm�+��"Bj�d�;�X���!v��>7~f(�kEV:K)���
��c�5M �9Rdv�� �z)��z�^�쎸zS�-��j�N��d�}N�M/�l��6�zo0��I�n��W�>א�ۋ�|g��� C�O�låD��>Q���{�W4�7B�� Eb��F*����Ы:��.���x
������͜�:�R��=�p�Wr8��,ԝ�_��jV9+·4��%�)��N)�`,�A���;��k�xY��%f������,�}u��O�;�cΔ ��F�K����o�C�N�T�K�}|S�vp+@!8GyS�@ce��9���1B=Io�U�-�KR~�xUJI=���19x�]�(?l�� �,P�lg�ʽc���Y��������{�.#BBY�5�u��nؾb�Bo��Y�:Riʈ7����u&��	����ϙŠ�i���|_aJ:�!������h#{v4�������c�|¯�O6��o���0"��}܏\|%$���8�G�`����q^W`�Z|�]K��\�L��h�7$p� `ut�r�9�GRL�)����j�����K���b]a�!�QK�u>#\�/�C����^M��	�C|�E7M�Ϣ�(FMEC�F�'��K�R�{&m�_~��.���Z��&c��pY��l��|/��Nc^�2�v�J��1N�C�����}�J�"��Y�c]�:et��Rwl9֡_���w�=�)�"<=~�� y�H=i�^"��|���Ið@H�ZC��®*���M��hw#遉�cR]'���&1���4,Ip#y@��s�Q�������� �����6�S��?Byv��GqY3����y�[���)���b+i�Jw�o��:`s3PL"�DB�1jy��b�`P��<nY�qsЧ�S�}ܧ�.~�c��<Z2���̘q+��t�lO염@%�cF�ej,�o�q_�)ĵU9����e�b�:���Y}�Y�ņ���ި!�|�zo���"P4��I��f�A������r��/B�֬��]�K+��W��Zშ���� ��k~-��)Z-�И�)�a�q��^�d�S&����Ѝk؉�E��tud�*�`���W�q�q;ټ���UR�g��|��dxl���5���R0��M�畟.�0)g��#Z�?	�:I7��U�h��=2�ݲ�R^�nCEzR�U�Y� Bp�4Dz�0մ�%�)ղ��އ����s��>{�K>9G�1Y"G&�}��ؐ(�<L�E�-m�e������Uɾg���"��`Y�,d=��c�h�ߑj� �kMFzO�JHqqM+���H��|�Z��Q�+�RZ�賵6��4��'�z^ȓ	�	^GB�a3K;��x���y�2�P{Kpc5�N-yVg�w�����U�$��] �P�K����CB={�֦�M}��r���dy9N�O���q�%����I����{�]V�9�ިF��?�C����bD�d���Xo&��[�s(��`�G�%�8��v�w(���ڿ�)2�x�9#(��"��xs	!�?Y���՚-����?͛8D�k���c:�g������l���Y׏ig�����JDR,�$�S�����-��Q� *��Q�4r�^�Zw)!1�rxq��K�<�O��"��X��gyXR��et;S 4WF���-���AR��s��ϣ1��=���.�l��}��5Z�%��c�"��L�Ñ���[�n�[`�;\����L�_�����`���!i4��ݼ��5a�)�d��BۄgJ�7��	��fx��߈��p��P�@�3Q��S��xԯw���(8
���YSX�J�.��)�-f5�����Ģ>�ջ��ŗ�J�`o��RAy-1��Ul�*���ۼ��%��#;�e	.��̣�ܠ���Т�-
�Դ����vHƄ�G�֌�	�k�-#]��]�4G�`������rh��O��P%?�ޠA�4�'�B�z���o2��ӥ�$����ǻBؚ�w�*�+�X�W"n8J��5�6�+�L����c��h�C���H��	r~5;�|Sa&x�%	e<��ٵ��Az���]�i�|Kc`�l�CW�20�$E�j��U8O����(�䚭�;���������Yŀ���7J�ޓp�Fwf�a�7S�a!{��-�;8�TFdD�|��Py�ز{����pę�q=�ep�_~8��G,���؃�RK�3�L�i�������|)c[`zC��l����!�I��V"�Z�StZ�+��/�N?
��5��fX�v�[�?i�G}���A�U'���ǀ/g��:<�B�K�Zd<E�ĶF�_yzV3�IId�X� ��k�v���!E�[�f,Q�s��<"M��k���LKE�p6P=1���_������7��)��^j=q呸�%��I*�ii���:ũ���A N�>�i��)��LM�a�|'By27���nϣ��6E;��� *��l-�������ܳ>/`Ɂ����ܛ�!�OW�(�W;K�4-�d�(hk�����������"�*۱��}����o�r�	��,�=�<���� ҔH��������y/���* �|�t��'p*ޯe�U��Ӏ~�n�{,���Ǜ.�t	�u&�RU�.�NoN���M��2k���]!�9�"��Z�Wӑ����D��$�o��W�EƀD5FҢP�k������Gl}��lI�?���q;���"?mʥUBƬ2;��3��ݢ�
��"c�n�?;�4� -W��ΣݖR�HSX9�}�c��-f�2r�a�~�rJi�"�&"C�-&&w`S��}H|�@u�+�3s�k�Z��(Oa^��SeU��>��E�X�]IZ=�@�8����s:T��2����I&����湩�3�1�mF��H�71�lbp
-�"!��#$��B8K.8��#!�U?�K��b� s�~J��F;h3'/��-y^>Ɋ-�ݳ�BM�欻�I1�)��z\���Nm���RQ��<Q��Z���"Vw�(M���䕨P��p1*I���ZtZ"�n9�\����@��/�5$��L��E���ȴ�ٳ$�\/:@*�װĩ�iT1@��҆�t}6e�$�3/塻%��)�����'1?K�g�KY�ZB7��:��L=����6���ﶅ��$���A��f�����u�u����\�	�XϹ��哣8��m�Gb��ɺ��N���K��ġ�:���6(̃+'��w46:G�2j*�s���$�3��'ͽ���1WU�����?����򒅞�����p�|D���M�v�c�ʨ�_����ǭ{�[�܇���pe�`.�j7*k�M-�ia �N}Ȟ��Iޖ�Q�s��D�9�2�W�G
�7D�t`o�Z{����٬��)��mG[�I���$�C�����a�S���M�*f���]p��� �Y���rY-o�{/��	:�1��i*$�=E�En�//	w�K�q�wy���8��f��
ܿd��+ɦ	X�S��E�ps������\���=�]8u6Q{��Vx�KIA.Q���i4/i�j!N�
�M���D7F�K�@�{������ۂ@w�W�Rm+� 5�#�J؂������B�֕�@���ܬ^��
�>�f�lE�����U޾ߎ]���z�p�'&ޒ�����Z�(��
����b��B�{4��M{c0уΉ�g8�Q �uZU�y�o��:�}ܾ������;˻O��;I����N%�s)��5���ģ�`�B������;�ݵ�M�X6 p��^<�[U����� ��j;��diT�)��ﰮ�:4AgH4k��S�[j8H2 �T:]���y�(�����pi�T�{Z4Jb����T6�a�3�U������A_T��R�����n:q}Tȍ-x�DhH�+��8"�Eq#D�=_�е�������ޔ�(��&h�3
_�� 
w���{���H�� N}���-�!�а&�G^�hݓ |Z9���cy|��cR�0����t.�Bꭜ�cG0���:'p�CïT��y�Ms1-��a^�k������|s�X>C�U����e�\%�=�c� �CK_�&�-��������<�s�m֪�=,�8~��e��ջ,3����#�y��%��%{�ݯb�<����d��t`���A��
Fl�E:t��A*1�2�G^�+cw~q��؜#��k���Iu�	(�s�e�����b�?]�k`��9歞/}�݃J&f��9na�� ������'������<d���K��Y��2��)R�2Y�;�˨��f��~k�]{g�r_~A4ǌ0�g �����N��@����I�,$��UZ�����:��<D{�TԐ8jiz���yğ�nbU��ǝC�.�V����zD�sGe/��H�����R���&i����4+Tߗ$�S�(ц�m'�\��x�ݎyngυ�gx"fQQ�#�g�X��>n�q� 9�87�������{�������A��@���Q��2�P �=�I���ߘ�+�нjS�7��5�(��g�B��'��/쉌�R�-r]�	P4��R�7���˴Vo\�ܓ�e5Sj7�a����V�qԌM�eI�hjk?���G�����Yi�k*��1O��UN@� 7�idL �wL�I�mx���d{g����*����)�*��_@)m���� +!�5�����J�Zuqd�m��f�~���ZY�0���9Kj��*K,Gu�n�!���@��������i>�[i!>Wz��}���넇���:Hܓ�~mh��9Gcts&�h)��VP���;_���P¨���p	XbƤ�x/_�5�i(v��[8��g�?����-�c;hR��'SՌ�l����{�����d�
�|1�XA����N,��X�������܈�q��p�e�)�N,��"K�8S�69G��*�"������6�~j�M�+�Y�e��m�Ah�"���- ��cމ���-sV/4���o}Uw��"��I4�B���Y�੽�S$����[����/�i��!$��߲7"�Sc�d� A�Ȅ�Ew��f�|ϞV�I�Ft���pc��1��zݮ�}�4�ncp�Vs�+J�9�h�strҨM����4���"�=�+�n� ����::1p��vS/Ul&�I��AJC=K��|���� YA�)R]����7�I����FW�x(���ZǄ51��B�Q���B�Ѱ�M"눂��X��ÿ�u�a�[Y���B��2oV��q:�+��t��/����i��FU�eT���L�������]ѐv��V���R��{���	X =�|&����B׷fâ������:H*�>�!��zm��kA�l������EY�sJ$�膹��o�P���?W��"��Q��>��󀟇�1�!Qp�1�gt�;2����Zz����H
�3nn�2���Mz�A�Qh�_L��BU��fn)Mn�
Li��0	`�dA	H���G��~�_�-`��} �ps��v��t��fG��Dx��O#j4��L]�ꤻz�Y{�ǳ&��4&sY�+\���k���\Xh�) �˘u��E� ��������5�֍�G�2u��$V���*N0���TQr:����(�/�3}��������b8}o�x7��'�_U�%�ҩ\7�I��w�57~��X��ݩ6H�E�ye[�!�}/}�s/\��_��&|�L�h���T�3}����WJ7
Սu'��r��~/���=1�B���ј�àw�ƾ_F��MV�����{9ё���q�=W�	[�����!��1��;0������U�"%�`�}�}�c�� }Nw�k�e�*y���2��>�%���LچK:��7`������vي?Ka -��χ$���;{,�woFښ#�d��+��g�>oN��S�
O�(�7#������g$Й�]A;����z�3KcF��-�b�m�0��|�.A邂�t�{ACӖ^��F��e�r����E�#���2mf���"W�1B؎�>j��0PP�>H�����|F�u^���Q�F�HuM�0O��������^��Xֱ ��S����=N`Vb!Wj��@�,2Ѝkrz����ڔ��*E;�3�*�9YcXՆ%'�=���P�ܬ��m��A[��:���G�Jb�4��F_��x�dۃ�����W�r��1�]a�j-v�������nP�o1J�ʒ��& =9-�+��I781q۵�r�h�.���3:O���לp�]�!'���M;-�f�= �9=�$+,R�_��q=Z���X�?�9=�L���k�l�( ����囑f�!za]|_'
%N������WV%ӿdb� ǫ�����@$+%��I�ѫbr���rz{d<Q���ʗˇ^��BM�h(*ĵ^�<�"}w�&�Bw�}��{P�hh�ꑁ���|��I�J�:�i��B;��.^�ֳ?��9�Z�I~�?
ц	$����L�:=�G���?vmZd[�M��MQ��X�w���D!���8��&+���d�We��w�,iJ�����GNl���QĨK ����ƞ���H%n-�3*8Oր|xC2^�����v�M�x�1b���2XG-�e]%N�7<�����)(j�i����U]f��9Pw�l���K����M}=k˹ao,"Z
�[�3kc{����Fuv'͈)����x؈93��PX���OPwv��9�#H���e(}j��b�6S�s�g��������q�o��_���1�ފ����ȕ��_����uv�ۭ������?�ڂ�W[h�}�u 79��	�e��6��EN�T����������"��������-/�t���`���e��-靨. ���i#��S�X��/�x~%��������>$���I��K�v��-�Z��n��<L]��U;�I{�C��*cX���`1� �r|���K�{�}Ʈfz?����}�u�˦��5�H��E�?��O��:���0r{5
�Yx��g*��Ms���R�fڴ�W�O�	�J��0m�'��]��x��
H��[<���sޔ��!�oؑ�@'�Y���E�bD;��`�_|��򜌛�A�,���
{g@� ��d�%E�7Cv��	yE����(vO�ߑV�/�;!���ҙ��ZR�nmO��6N1o�,���*�p�����Y?{�؛��z�N���$��0:��@�a-���?���sD̡��m����K})�U�>���r�DQn ��sr����:S���x�zF�;�`?
�T��Œ�����4����wl�)���
V����g�頪�J��w,��
ׄ�Y�mF�KqzA�j�W!`8^nf�	�*�}�ש
�K������f!@��#��w['���T�?�<z��sן����"�O�8c�u-�@��2�SN(6�C����(��q��+rQ �$vLM:3���N�F1
&
�ERX���=�!���L昬g���H���h����:��8����^�|�-��r���Op�5�!(�$�:��I~,��%Wf�Q�;��ϯ�sh����=3Ý �![���-��v��W�L$ڞP��W��r[~o̕����N1�j����z)�@��s+>c+FZ[�']
�D�@�K)�!���}�!�<)�˓a�}����V�A
#�Ԗ��(�BP�N�ؼj����H奠u�f��}]��m��0��Ǵ�^��BvB�Wă�(Wj�?q�v'�i���[AMcQ�����6�7	��*����I���u��v3�6r��b�~,1y*z�U'ә�שE����?�T�RK�ɳA
����xl��P)�.����Ѯ�����'��ͱ��Ox�~�>G�8�?�p����pd|3w�t��]�ѩ�{�������4ܐ����M`غ���S�9I�-�R_�bH�:]z�ڬa	�S>�3!�n� �����n<7 �.<�I��^��Bc|CI��xvN��k��D`��f�^�pA83�5=s=�O��ڻ�`H~P�j��N��u�F� O�Ѩ���6,�T h!ʨ�q���p<'F�%�[ހjͽ��Y
#��ɘ�R*�6���%�m/L�;�F�0,��}��~��h��R{9*�Yd��q 0m`g�(����������@��������p`���nv�T�qKA� �3�d�2�Q�5�i!����
I���KҌ�0/�4�"#�$���[��u�W�w+��֞�@M�>��~~��ub 0U�tMpZ�i�m=���o��5�~z��v�u�����["�c�V��(��9]���*8S�Է]g�����l҇/�:�̨�j��mW Q-��"A��#��W�=����Z��#�M�t: �e���m�	>,
]�U%����o�m�e�����x_ԛ��O����ba�����%]��z��jئ4���q-4b��m���k������W�0��;��@:ss⤝�?ف���c;P�H4E�ZdBQ��?7��7�TV�4�|4?.�ׁ����۟�$ͼtƦ��P����1�̹
��|���N�^�:��A2�"4�^�}Y�!	��>₊�{S�h�Oex���NU�%W�'1R���.6��0|�p���V7�t:���r���!t��VV�]����?�Y�k$���v�9�^��v��8�;k�8Y� ��$O�����,Mj<���4�)j;mޖ���/���g��IPx������_���xO:��*�5����KE| M�b!�ؙN�sH�❞�'�٭_lS`�%MMnR�eoi�/�5��϶y�T�!�ÿʽ��Ż����&���c��6��/:\h��A$&�RI��il������J��]��!-�!PCd��}�,�H�����V�>J����Q�""g�e�\����<a2�\��Ȕ�`��s����LL~��d�`�
���8�&�?yiN�ǽ+��N�@������eb�c�}h��iTM�$&f�ox�&�7���Zuz��8N�A"���Φ�q�됍�1�)	�PX�ϙx\�e]jE�P+�u�ۜ��VzF�R=-uBO�PQd~m
$�J)Z��NW��s:u�٤&��Ey��E=���.|1R�	G$�6z�8 , ���9������$\�����ıI���2ΐ��~*�O�f���*Y��_Y�=�!�/�q`����;� �JII����;;��t��Mh��6�Yv�Jg9i$�F"`]"��Ys<�3��ӯԀ�-�95SBl�>��ðF�'����7�35!�P�[z2��K�"��߮��yݤV�g�[����
�3�\~T�=ש��P��SlE���g6p(��!2fZg��p.?m*���92f�/�q{F�:1	�X`X-�*֎"$
g��v��C�7����F�@;��qx ͯ��f�k;K�I2)�?.��%L%X�'�یȑ9+�B1�>�h��2l(�����ǅނ	��`H}åAmp@�\�l�3p  �����}3_^���PN��P��"����_�2���fh"��w�JȮ��J�S-]�1�j���p�A�NF�V]Bh��&NCv�41 ����唀���͏�s����\5�7��f��ͻ���dU�u�C�~}Fꠧ I�W�S��Pc�߫S��:M��F3���5rև�����ȢT��F�ɞ��ecf�=v�Ǐ,�)j���6��z��C��BcCo)P��m`�Q�|���aݛg��	��U�P���̩
�e�<oXe��>�����}�%��qK���3^��C)���h������ѝ�6K�c���D5�ޅ'&�Ի�ٙ�4�����;�� ,���^���x�����y}SūF��N��'6�څ�W!ŉ��Z��I�;8a@�t�x{J���r�dJ��3��
di�삭�E�t!H;��.���t�%�ͳ"�l!ʱ�(�:�K��L|J���p�� i*��!3���, �fB#�����AA��h\P��(xz
)z��HK�&�;������.Y3Y��{�(�J���P	�A��N�XI� x��ψ�U|��� 1�gC��h�L�9'���]�K]��p�cG�+n!�Q�e�c夑��z]�چ�ƝA+�f�L5�,⇁!�!��������/z�-�׳1�@�\I���"��C�ߞ�y�r�,
`kNA� x\�� �N� ��V(E��ќ�ΑF5�0yS�X+*[��#�B�6 ?�y��s��xtjX�~R����i-U=�^W��B�_�B�bm'�`s�bWRUpi#Q��-ur��t�֩`.ck��C�<���4U�JxQ�&���
ʝOZ�(�s.Ѵzp���R��JP�J
�qK�����o�c2���>�����1}�7������#&e�T4v̈����QP�ؒař���2]��{?��tP/��Nv��\�\��dF�2ݦn��J�qp��^yk�L<ʹ��o���9��4��37��5H�7��5䃖���<��uSʔ���BbǗ��\,NoS�H�J��#R��ǆk���}$��w0��Fk���w�2�&��,\1Ϡ��ݍk�>��]%�Q�y����&H���i�E(=� �K��������ٿ���	Z~�K�Hܑ��f�{ 
�DOn6�����ם*�3�lJ��xs(����}]���_8�[��ܔ�&�6������J�}��o������L�H�~	.W��$�S�	.1,�VMalJ��L����L͸MGϑ����n�-��:+�S1���(#f]����Ij�O���il�	�&�b�~P�W� D��s�P	�F�^0���f�0a|R�i8.u�=����p{�a�3}�,W�'��I�f��vd��13!()n[�\Sh DM�R� �/_D�����_��OC���﫭���g|?�Y�K߸����A P��9�B��_u�8"se�c�2�.:&f��� ש���R/��>�=E���1������ӣ������XG�x�(�V��z��1>��m�'XW_�ꤪ��MZ-�+p���9�����Y��ڇ����`�*<]z����� ��&%g
�-�i��>�#��Թ~3�A�P�.snd_3u�J����H+k��&�Uq��%�G��G �����3`���H�Ip׋�̙!vDî.k4+F��e���r���'�W�D�\3`�i02���+��Ś�zLS�6��m�0�,b��dE�]���LY O��mF����*b �	6I��p8=M��m�PJod���4e<�o.��tV�yx��9R-�����{����ʝMiJ����7d�V�3!��|�w){ĨJ:��'F����Q�LX��MrTw�!1h$+�'�|ư��P�8�0Q15���I���,aI��2V,4�v�Ѝ���(2h�b�{�`�X�S�*%p��q�.Vl&�o#;/�b�2��_�LZ5�=�����1���
���eƣ5�j�,��;݁�-��A��cMbt��e�L��6��QĻ�\��r�z��|�O����Ga��ȩ����-N
4��Ny Su��K�aJ��B���������K�uV4
�k�=۶)R@E.%��i�u�������f��{�K��x��R�A<�jΤᳮ�L="ȿ�%8F|w�Q�q����� [.�r �hq�O�uEa?�P��Ƴ�����T�2?�0$?db���#��>���+���'�S�<����/���=3�������*�#p�|�`ҕw .n�O(�n��߇�v�������"���ߒ��'�݃ �+��R ��6C�c��#�����  ��Y�W���g�]㨊�y��Eg����!���ꜘ��ۧ��Ks�&!� :��o�U�ֳPO���.*eMB�����8�>_t蘟N�s����YuA��M����xWU��͌�}� ��(Ye�?)�%Y����XӰ�fg�9�ٽ�\|G��MF���e����J�~�Gശ/�Q�̽�)��� Y켱�w&���"!N����.�ĢD�yZ�������Fg�
=&��
�d��p��w�%�r��(���K<o0/��Ӳ,�0��$����XE�Ϯ�4o`���ܸu�_Q���P)||�q|����
	!#&�U���)$�~R++&��Sb��)�B�����ە3�_<��,ܫ��LrbT�鬣��p[�o{����7&UE��.��<p�yO݋�������ݷ���r�l;%J�I�h�R
Ҕ�Ę���ZD��c���*��r�/6{�Qj�{�L��pP9�p����ҭ��KP1� �g�[�����{�j42+���P�YSE��M#-πCs�A�oÅ./f5C'�P���r'&�4@�-���}@��'�0ʱKP%���N8e��f�V�oLA���:�U.g���_�`o�	r6KC�Bi�5o_�.�a!�A�T�����K-e?<�qL
���~^�aQ���Gi�^��	p��(�g��[���Hb���҅�㾽>QX�~J�ÃU���*��93�`*5�Ȯ����a�����MY�b#_ZS|o�o���n2����d8��'�jށ�vS��k0�7�c�S��Kv/�����gO{\�L��������ZU欄�-����2:�Tp�Z.9�زaf���AJ�^tEo�0�:���P���`��}�tj­�3�=���S�4MH�^J�u�gŃ7��;��h
k+ի��M� ����I
8�����24�G*�2[�3��;����&|����r�3�N�)�v˽�.D�_&m��X4��7Ψ���L�ź��'�����|1�կ���`��	��
i�l�F
����+�x��+Dj(�LU!
��҄�#�s�.-��X޿v�#vl[�'�$�M������C[��l5�<����-���Dj1�yY�w��~3�`�	��,B?�[=��B�R���{��g�Q��jMb�\`��H�D�Jr	�8�g����qv��d�[�R��?��h�/Ǉ����G�h��˯!�iNe
�s@�N�-K{���3&Mt}�br�L1���gp+�+tc
Y�k�4Um�����Ց6f](L��
ƒiFګ&�8�/��o���4A��T�����F�Jv,��ӎ��j�j6]u��EPz���h{#���K���0>���	6t����U>�'�F:���
'ܢ���%9<�n�����u��EM<�HJreՄ�il����C��[������K(�bN+zys�V��a gQ?��"�y#����Z�q�9�Oe��P|k�e0���P��Ɖ�)ՠ�����3��#ʣ���Y���	H�~�-��EK�	h�w�����#�S�;��zt�l鲕"H�b�<�u1��<Z��*$���j��LMo5E�������&Ya����8w"X\���L`QT�q9>�$2���{����D�"hO��Ff�ō@��J�Q�`n�>�����N��ik��K�V	C��W1Ra&�,P
%;���G9C�5��P ���pə�葨�l���C;�_
C������� �,�x�ߨS��c�'_�� �;��dȓkh�M=0q�S·����/�_5����5�Z� Q�^��rv��8���Z��s0MbA���= +/�T��ON�4�b�� o�� �d�N�����v��Z$�Z��e�H�3Od}�8ڡN�b�k����A�Q�Hi�N��=&����
�Q㞹�oFKe��n��+��s�%�Vމ�Q84�'��I:[�rrkSfȀg����u�7�at��c��eB�����.]ʥ[-Up�~�־+�W4fD�U���*�%�yC ��/�Rmr�1�/����6i�fU���8���;Ci&����T��y"*�*/�N�A:�GW�e�g���ȷ�E�1q*P�$BqY�&	���y��8�k���-#(7���Q~(G��]��Z�i�*0������ɱ�$?�����s��K�0Z��㢩���	d��z��
�VlHuM"�Ü�Ђ���A���$n���^a�S�d_�����j��!_	��=�m������N}�k���C
���rva����g'H&-�fK+��.�A	��p=Y|�n^T?|��kŸ[��S���!6��A�n�s\�զP��6Ō�^������������p�%思�c�Z�h���+>��v�0��q}MT7ek���+{c.��W<�j��t1�XTe�?�U�O�7,�I��.�b����Qo8���������]��7���va�U�������%�V��l��<��L��,<�@i��|�K����~��rp||7�����0�%�}�=�qI9��H�X�d��T"%Fm�|�X��a�x�DjAz��[�����ڶ�X~��я��Vw&�z��m��0T��L��l�E~�݉�z�z�]@��&7�#7��+A@�a�Ns?��!@�[ r
C�9=4Ć�X~��A{�ep@�ޓ�v%[�hL���8u��ڤ��vsL8k���>�����l�M�����]�GK��9N D�49��s��WN�|�q��PoSg����(���.����ЗG��M(����L��G��m�z�IM���!ҁ���w,�T������M�3�l|�/~���@�j�=��w�^���ӜS��oϑV��PP��QM&e2�
�&\��i�i�������2�	�Q���s���Q���&Iѻ�����������]����7�EZ��mtz�HHl�+V�� }����y�R�k��Jba�*�6V��Z-b�<��^-E�f.]e���b7'���q�=�!� ��x��Se�W����c#XΟ�o�\�i���Gc������U|/�G%e]�I$�џg����i�����y�*/��!�z߄4أ�����L��<�G�ҍ#*;7Źr��vڹ��㹰�dM�� ��P�(_<�@�ǯ�5r��k�����gg�O��:p%@���ZX�=T[�5�"蕈0?���Ml���S�����j�u�KV�&ߌ~��@�d��?�Zf}��o�M���W�_sBa�b����w���b�yd�_���P�K#?�F���-�)b:�"z��y��Θlg���g �oY�H�[�E�$���h��B�.<�	�U� Q����|��%���֮�c�����w�P��	�9��M4p���%���*��|vB��@g&vj��n���MN5��/eu�r��G��h�3K��2�s~��N�H�4)Չn)�<խ=�s4A�2 ���q������
�FI.��4Q'8���F�w�{9ÜI��¹��}΅���*}�wUv�}��"g-	��%��,Z�u��֏�V�0�z_�^��(T������|��3B�%��ض��H� �P�����o[�~7_�~2ML��E����%��R���(P�CA�4�#3h-}���T-J��jc6l�zt�,�x���Co���7z-��T^MỤ]	���� ���/kV|�Lq���c���6 �ĿA��Ѱ��Όt�����{���X"��6�C��d���uVC�u�7�7O�6_�����%#��P]eg1iC�Ł���E��+1�V�@.�x+�ڍ�>%;�ޭ���'�9����@?�N-����N�i	��v�
�䝽{m%���b���&���-HO?����Bd�� ��c1o.iC"��ϵ�ƌ�M�
�e�i�s��H'4ö柉#Jx�ۢ%c�$��#����/0�������ʙ\�*��f��=%�*#��'z�R���x�M��3L��!��0�^7��~ۨn]�)�F�����um�ʘO�����!fbt���#櫋��B]�K����zJX����,�L���ݢxfE�A���짬�+��F2��Fc�/x@=�o�[V^�Z���OZ����Ś�YU��Al1r�7����e�V���n(G:�Ь�L�>dt��m5g֒��#�$O@�_�� ��rGD���6\�ˮ�8C�2y����qh�c����́���Y�l��(\}�Srw�^`lH@=�*�w&f��9��j�W�/cXp���p!<��3����f9��?t�=I��oV��٠O�ۆRx7z ��V<�˜)R3�t��i(�r�9x�U ��-�8B	2��l�8�17F������۴�A���HOx�5zywB�oR�x%�b�s$]/����+X��y�@��Y޾�r�[AK �-� E�!�����ZQ���Gb��������x�K��#L�_��O��dD�ީ�Ja�@���,O�q�\��49Ol`�C��y�⥽y�Uu�-]�Z!�g����õ�H�uO�\�ڲ����LJ�����9=5�<��{��y1o���2}�nU���Fů-}����tܬXJ�p/�`�}��{�E��n�4��� @�c�� � ���4���m�C�_��}r?��A�FY���H:��K�aE�z�!V���G����c�Vr����/��|�طs�u#���DU"�J(*��}cU�J��D`y xm�m�F����Q"��^�w�]��c���\Q.eY��T��k	-��K9�P�R�P�x󒾲\���~cx�i���FVǸܙ6��b��AwOg����h
�E�!,X�V�a�"�DOm �.���I������,W�.�B�~��4�fAt����֜FdE4���ߠY:���d�d�M)&��}Rs-N�q"�\��kڥ�,El�n��6u����2�4A�У�����,D8b��0�B�'o��}q�j-6ܻ�\��nL���q+�]�*z�
?�O�N��lG�x|�p}6�9��	�2B]g� Y��5��u���'I���yJ�t���v���3Z�^Z���ЫZݝ���P������{�o9)�'/6ׇ���Y��rR,a;��j_��U�̢e�E��'m���E�[4t�S$�1V�1�G���-�:e�Fm��P����rhtb��^\^\�	/�
��Y�K'�G��"����L��i[A��Vq A}�m�Ln��Ծmx��V`�u�*���ͱH�+[r�fO�x��?(V>����Qڹ��?o�G_?�HE�I�wQ��I)u��Wt��+e�K������l@��۠��l�΍8�ک���!m����v�6��$�d^���&18�.y�H�u�g���M�*�5i#H�z��2ƞ�?�&���v_��o<�3wo��c���b�1��M��!9�@��>9���-9w��l��sm
�#E��]��v �����y�@k"�G�����k������L��ϖ�ŰMYP�΂��px8��u�Qsܘ��4P(ҋy1*2@����O���+R���+h{s4�����π�D������@�p����񄑰���)��jCek��C���� z��=]��X�MiU�6x~h�6�M40��"lO���*����碻[;�X���P����1�e��X&�(x|��]��"�Ǟ�	��ʙJ@���'vI�/ň-n�ޒ5���:m�SY���O���ApDկ�O6
�V8��`a���i�u$$
(3œ����Z5�pa��ƺ~3�0�Q
����I	�e��!�S����������Dv��t	sAj�9���#C����uD��
t�1%�/���\I����	�<��`�X����Hػ��#�z�ݽxp����oauA�W
ÇK8�³>�o��j�9v�b��,��xQ于������^���@O���Vㅇ���+��ֱDdͬ�����3ݪ6��'���K}Ţ���
~����F���CZ˷쁹c�[E�1j���{���[�O�/���ob�<���~���D�Y��}1�?f�����3�|W%�$�}jG�2r�E��[�ng�˞f�Cv�qz`�
�*)������_wZ�k;��%�`��d��B�EK�]s���&�Be�(?i��|�O!�.�F����X\��{[�~�N���K ���
��E1��b�����&t��X�5�q�/V��wm��3��=�L12bf�C��*WԦ�; ��5�V�:�z� ���Q�ݬ��~��ƚp��*af=���f6����D�,rN�0�����i�,�``D�bF������k�<4B�=b?	�3�e�I�Ќ�9���`�_��w��r_���T\�l�=,�1P�ҷE����ݯ�z�{�ko��p�}�h��#�%AllU�I��|�Hk5�FA�­�ab�/'q�{��*�l����X�XG���=�FT��"L�g�3D� }���n��`z�Y8.V�X2i:�7���!	}Z��I�U�am�����]�ZO��_!��I��H��E��F�軽cԀ�rH��r�1l!�����f�4[����
l��z>1�`J��w��,Ƒ@�8�aLx!��%��R^��yPzY�(��,6�e��~�C�tad%1Z��O�ܵ�ʔG��[Gb�z�GK�>�h?��"�),pL��y�� ���b�{t�~@����jdH�P]��1RSJ�&�&a�	[�U��|	/�Y�"���o������(����*|;���F�Q��U+�S���'�C���v����#�4Ȼ��ŔZ�
��\*f��w��`i��<��'��g\#P
?4q� �l,�+�Y:"90;�.ٔ�C�_�e荆�8��t�_��l:����l�����|���� ~.��	Ch����4Y�����ؤ$=��N{�v��H.D�)�ն�/g�MƐuA����i	r~�獣K�?�c\u��-[��̨�.�;�ȎG��xN}�;�s6�A�*"�Y����Sim�OX!H{	E|�D~3ij�P�-MƭX�\Q���������h҅��7
��1e05("�Ŀ��!Y����&Φ��������t;k�ng�I�)c����Umj���À�>dܴ�	k�Z��,��B��YB��f#@���3
�8�*aݹ��:,{rw��e��y�H�q��q���z�䢁*)"9���8�`O��T\���g6 7#�Ũp�O�"�Wd" ��@9*}U�		�0gđe�DzBjoON�	]{eny�,��l���
�C��I��No��7�U��o��죕\7���S���j�_��#/*>��ɗ8�DD�C�1��ɖ�tR�gP�l�rê���F�*I��u{U��N85I$�m�F���ۜ�,�N�D�V�p��L�|=�\�1f�K&;���ń��dR�a�s���6J��g����I�s,\���N�YŬ~T�7�������R34��̙�7�µ�	h����c����wxC�v�z�A���<JBR7�C� +muʑ��=���~�կ�N�z�O��՚�!
l���X�'rW�TZַ��hw�������/��E@�)JX�9x� �t�	ӨC�^���8�
b��9ܠ�}�]�
�u�I�J�H�p�?���7G�Z`X���B��m@{��A�`����*��9S�OJ�+L���{�T��M��
�	�n���AleN�`p��]��D�LJ&O�J N~� 'YR�ƺ?~@�j*�[�t���t`A{}�<E��k�҈�n���V����w}��>��Q\��,i��m�Ú�B��o7
V7��H�9�X�0��s���U�,�6�5"�3�eKHm_Y[�^x%�ɩ���I�6�e˩��Ν������$a�U@4��ͷ������wM�	m�kB��x�YʗE#�X�섖e3�!�-��?��J&�'$G!�}֑&n�ʞŔUDFS�Fi�#��<���	�^7΍��&T�1� VpZ%��o��#��x~9�.�>�_Q�8�����@W*��E����)V�S�Pj���*b���j�<
y-�'�6j�?���6�x�rB�At��ډN6肇�in%`�I�
)FĘ~e�z���+��4�sD?�#;\=�H�5��G��B%�9�C���@G-£�W�E%U@4N��� ��#�����T�@�x�����m��LK+���@Q��TO�b�+ƈ�teE��A*���kxk3�J���
c��"�7fO������A}m��N�0��3kd��gZL�N�>Z���\���TE�Tq��Ң?0�$HLE�T��G����D�^m�Xʯ����(xjB�N�1=B::����8�"g'�_u
�I�����|�����ˢ�t9��Z�I�����R�D����0�
x�bR+5�]�sF7z���/kF���e�;�m2�kX�t����d6�	/�I�b��p+�F3M��_�F�]B����T�ב&i��Kb�/䄜�_��Iq�Bk�_���+[��`3���$l����'�����H�	�2�A�����SH�v=��/��:C�.�0l��DK>K<U:�ș�蜾��Շ�����מ���<isR;<P%iz��w�U�XuP߸�-�s�d��ԛr�5}&u�qL�,�o��9��k#Ggz|l��9���]4U��W,����H,!� 'Y�Z��N9��Sw�~�<:�Z�0�����p�5��uzyGزOwҶ�{�1��2|�5��$\kb�t��6_���j���9��Ygb`�#�4����v����2����㸻uy}�����'$=h�+D~���/�y���YoF����07���Y|5�,��=��[c _|���Vq���;�$��NlKj����dt-.���go���.Q�����`�V�=��O;��b��)�G�o������x?̣��P��@�PŮY��N�ib��	�p��Qѕ�R��䈩Y�g� ��2M|��륺V���t���~�<��hJ�Aq����x�����j�U�\��8H���8���3N��H>~Y}�L+-;%D�~��.�?�BR|��>e'�������Υ���" �A�Ϭa��>;;�x��Mt�)����/T����D�~�J|�b�u%�����^ۅ��?�n���vlO�7��_$U�GE|\�4]�X\�Ԯ-'Q#ՠ�ؚB���!e������I�DN�A���I)-�!����;j�
ɱ���Tv���^��u�xy A-By0
Q����2!����1�v<�u��o�{e<}	)�S����v��j�镝����3m��-�� ��Z)og	�0����E�!��y�b!���܏��v�S�������y���t��7$ËZ��(<}��� 4�AWkDr3�����Y�Q�:;����!^ˆ�e�_�D�7�CA�KӤ:�h}ڴ�`�$�L���4��or��[��/��dNR9�Ru�{��q+f|�H�V�I�0�=��
������Q�c�Cݶǔ1��奷C��j,(�م LU+�?�J�?IV��LP1������ �z�;��
V�4uv����}?Qc�:U� 2��ڥ�#.��_ o*��mK$�N<�}����h��/�i|��EL=��G �N�[6�e#9�U��# �ɜ.�q�N3���������	ݾ�p�I�3����ʯ���<��7;<��g�ԾX7ْ�6�e����5���͹8 ��R,��G���	����󜷵	�\&�� �s���,��Σ����C���,=�\k��{>&�Z�̬�Z��b��.ǎ���<��ܘ%���Km6��`7d�d�%oH'J���a�a�K�#���f�L�pF@��'#|�e	A��K��÷ԋIf��#g�a@s*�{��3�M5ut��#�`�o���kƒ#��
��ʐ`�Cb���A�^��[��Ɣ��|v0�l_C2�ה;�I>� �9$ߡ�i�q��ʔBl+���J�����e�<
v�ɐ��¼m��1s�	�����Nd4ڸ���~���Qe_�vnJ+��j����Ϋ�����R%f������V8Uy��>8AO�W�`)�lb]ж"N�y@ �v��-(�囈82�X�<�O3w=8�0Q�µ��V�)X���[p�o��/o��7�SP4d�@ѵ|�n=���Y��
��K��A
�z��Ϥ,�(����x}<��9RV2`�k�Q	�a C9�����fʪ�����d���ÕJ�I��h�D�H��>���s���8��Z�U���0H�[�� �������諟�B��V�e���@���~�H ����ʠB�-�X<��鷹���oѭ�j��z��<K�����%��j��H���?6wp��c��"���p�Q�T]���m�;c�����������i����k�I;c(p(_�Ts�&�M�<S8a+�cC�9H���a�&�%�̎@0��L�O�)�p~1��$���	{/k7�<"&�$PO,иkyS�~�,9!����g[�醴�HA�kl�G��V�E;�0p�&�r E��<��B���EڠK�cCO�/AP���#_?�Ⱥ��đ��N^�t[l��Rn�nY&ir�[�k���_��o?}�H��(����M!���d�R˼Ji� y>�?5�B`���3TG�����\�ÿ._����V����#	a�5�z'-��*hf�E���݂י�B��"�4�}Nq����1gd������IĤ%�R�J���(���B|4k]m����|��;���-eX�q���3�y���XLx�#\О�V��d=���%������ �ɤ=H��)^Q�fۂ�kBe��>�Q�)B:>N�����j��J�+��G��e7#��g'd��+60�;lS3��m� :���2�xm�Z'<;~:+�'p?ֺ���R�06��R�΁e�e�KB�d6����͑n`��"*S��Q�W�G<_I�;����cNVMoo�@�;e��%jv���g�{��d�L���y�5z��|����M0���b��j@������8�T��h�_M\�S�h)��CWD�Y����s�1���On�;l'���ip���>���u^��z2J��E������΄P-���DY ۶��Z��␵�U�{k.��I�hw�N��n�������A L����B���7wx�!.�xI>�؁7E�%�͝��z�x�'��zN{�#�u�V��0�n�go*[�Wfc.2�I�9w.��2r��ۑ��s�͓QDf�˭�p���`���� u�//8�uw	;P6�"�Լ� .���{�3~MO�X�Q������''-N�,ߔ^L2ǭ�w7��Y���E`�>t�����~>f\�g�>�'�UZT3ir�W��s��x*�^J����05H�W��L�A��h�;&��w�-�/�J�T����-�D�Z�9M�������K����*o���0����r��"���Y9945ѽ�����R��a�X����Vf��?��B+8}�?}��?�qv/KE墣f+ڈS�p���q�
���Ł���
V�Ga�;�i�M�n�û��"޾w���R��S�r闘2o(t3?�o��lR�]*�n�fhQ���@����3��OW]����2���N�)��Aq!��+5o�[!���w�{��K�1(��<���^���c��?{�mh��[u�?��P�Մ�Vj��𨗭 ;��Mg\#m�X�>%��
f�5]`Pexm�,B����V�nK�j/�=�ٖh�&�}�Xe�E���2�*/�k�qt4�%3R���aκMW x��z���  	���	(�Ț�:���a�0OƔ�/�p,t��/����Ձ�ɋ�_��������I
�\�Z���a��N�~tJ�bgs�������U�,A�#�9�j8� ��!]"[�T�fgeM�"T��c�,�����h�0�пRu
��S����x�Hf�9�jk���MFUa�6f!��
H{��E�0f�ge�p�����'pФ��4.���H��N?<iP��vx��;��!lB�'o� ��L��3�_��S��V	�_^�Kί?��H�06�6�M���x���"ێ7�*������Bߊ'���(�L���� p|\��Fݜ/�|f�����4WS C�+�������צB�G٪�O�ՠP�e�{��A����������j$u'lG`h�����jZ���C\OZ����� c򝛄I� ��U�p��3�	/�-�y ��D�!p�*�[Gn�Ȉ/�^������/����yX�������°d7��d8jH�� ~{8: ����W��;�YV���8�t_o9�m�;ػ6t��aY�����6��T �#�&��u�2â����p�y�ͣ����ֹ�yCN�z<^|�r�,�u�G���>u.���:��l�KT�R�ڝݍ*���{�m:'U?+M�%B��:d�b"4���P�95CLs��Z��mw@��/�H�2�HnK8Q�,�я�*��NzL��O ��P�Onq�]�]�o���H3�`�׭�*�Z�u��:a��R����<dS��H�\�V���$[��\"?���ѐ����
uG񡤨ղ�_�O��Y�0�I���'4�����ڌ[!�Xߔǵ[��YS�o�QGN����ٌ�<E�<N��q�n>�E�n- �5�0�RU��"� �e7P�"����*���U2����q[��7�4'��7��[#o#�e#�����E��E�6����~о�Ս}����.�-�A�@�����] ��N�Rp�&��j&�(8�3�[�_g��>�f v�?W�-��T�R�U����uԃʆy ���A܍%Mc͏�<:��/ݾ�u��1����4�pXH!%T�&�&���٢�݊�hS�B�m��qG{����-�;y�!t*XS9�c�Vz��
I�B?Æ�ԗ#�j������g
%�*�O$� ��k������m�?�_]�R�gYF��lx�扙+�	==�K��8I�k����qDU�]R-u�e��C�+*	�*��+�:h�])�r��z�m��>�lP;I�'��>��͉�ֈ������S�'#�j��~:�4�xcj�)e�-�$5��џ��]hO��)�r�����V�hZ�����c$Z[���C��RZ��b���/��J���Ґ�!d����n��5�Cuv���m�5���|ӻMG��k>�TȐ�K��ET���$����e��;��Ё��D.j%��/y���̋m�O��T*���:��:3J;Jܨ�t� �'k^��b}Q�8-�w�ޫF���Ǉo��<��<|�vm����
����9���b;ō��g�J��/\���F	.��w(�����]�N�=aL�~�Ü5ajQ�k���I&}��-n{~J����c�M�z��h6�#���|v��O)�u`��O��-)-(�."%-#Y'jʘE��@V�k�t�"��NI�K�t��b�����a;?�:v>���c0'�x�j�Y�0���X��l�Ʒļ)i�M�Ag�# �3[ds�j5��=F��.,�����(�D�Z���b�0�j�]�k����
Kn�`�7ujT��z��%��Xp�|L�SҟI�~`Y�_d�SQ(Gȑ�4�B�4I���R��26dcwG��r��i��<ƹ�^���䣕��q�|.�C�0d\�Jg#�ӛ.��gn@�	�!i��j�C�=�XA~wzz��K�R�*=�=�T��w�-�*�N�Rpρ.�A�n��}�o]�v3Y�K~Y�؁�d�ZG���<gfaĺKB�:l~�y�J*�Q�B��Z��O���g톊V�����l�M��_�=M(�棸�{�f���c�05�㝏���	���Q���bn��:0HU��raҾ[�Cy=!=�h��VDʬޑVKh�_�	$��1��$ߕh����~,;���lyF#m���p\M8�[�����Iז(��s�<9�Lv:1��F:Q�@�O�|���8�k�����Z� %1����e����,�	�C�@��BƵ%!�C/��S�`����[�6^�;��7B)f:��9����K��]��m�A�N�7"��9M���$��_��*��N}�=�{?��J���F�:�}�U	I�
T�Wb/çD���r�RՌ:Δ�%�1���{O4�)�8�O�,�s���_:=�j��)�h��94Э������F����m�Y���J�φ	y��$x����ဤq��|��aG2���J4@����+3��mN��#-���ŒuK��S�����mnǏ�-d�Q���<�i���C!��xhH�bN�A�xY��5Y���8^��?�����[WH�L�{�� ?�$#�����x�ɩy�h� ic���E���5��j�B�D���R�j�$T���S��U?Ί�%aS_�}�����z���v��c#^���u�6���ez�H��tƃ}]~��0H���b�������Ή���׸d�#��������3�z�����=��h>[��(��>)�� ��f:��J���m2��z1�'�6�fn)7t�E3pj*ۻ�����s�<P`�tn��@� �y�g&�S����W�����`"1� 	�Ǣ���
�V2�	m=an{�����?�旑��䤑+	BM\�?����.6��sAnM)�wM�e�`�$fM����7rZz�5զ~x� eu��TRo��q�%$@^2A;B�*���V��*�������4"$uD�D8��&�4�Y��<>�:愑���#�������B���wyߴٝ����Yp��%���ܰf��?ϛi�|�DƕK�� EJӐA��-F�u`�]�����W/�Gϕ�mEݐۤ��Ŝ`e�z�,8�2 ��+=WI��NU��fS'��<vz�t:ge�v��s�6F���+[s�
G(����F`����}d�S����M�>UT�<5��m˘�Zr���i�'����n�4�A����P���-jM�`_��!
)|~�>��{*Z�q�)N�,v�y1�;��*/F�$�c�a�ZE�Ѷ�4��9߃���QQv�e����A{6���Iapa�7�� 	5��LQ��RC7�7�)?�ǹ�T�xFc�떍+q�k:����5� @���5��)�$�1 �c��=E)ԡ蝋vD��GΩ�<�8��-��+��c��x^�Ko�3_0I�d2q�.MS�F�8!��C#�g�`��Y���s懂��BK�J�]m�,�sR]��44�dU4B��g<&*��+[��$�o��N��XEB��&sң�{�ꡖ,����J=�_��n3,��Ĵ�I}�&�Y��*��H���/z�zi�6�|g�֋-�2��ن��g����z6�5r�\N��t���@�"-5(D*�˿�$#I	N}��_ͬ'd�6��4e���s��L�o��]E|c�I�B�x�2��"+���N�e�@(_�7q2%9���s�?RWH�M� J�����z�I[��0 �6d�%�ŲG�鄑u�%H7t���PE�`���a�rڽ�����l��$1oU`�9���$��i�i�[��ZJ��)�д�S�S���*X�
��=#J�Z(����X<.�����
S��y��y�'��� �x:�=hfqתaOq���b��bl�K��@��"�TKE� 2���9���}(�L�3�B9x���S�78�"�*�F;�H�kq=��/�L�����-�<M2?��Nr~��%
����
O�����X����~06d\W��%5l ��;:c!S ,'��ρ6k�i���-ՠX�kX�R�E��E�.�͸�vˤ"%�q��l��phw�֜�.9+�'�o߬�;��L�
��-��Av�TN�05581���bA������We�k��4�W�<�C�#�ڷ�?���6�[FS��_P�5i`?n��7���eK�y~�dTZ���/&i��d;��]9~�%���熵���,j���%�*�*�ަ8�NrL0���b���%q�
l��/O[��i����2���O���-�ʑ3�|I��Vk+�kJd7/����P��8��q#{@�i�@%b��?� ^���/o���u��jߞ�),��|�Y�r��g��%��ً���{��A�_�T}���A�=A��8���Qn�Ŭ�L�]~�A4m��$g�2O�mP9�R�&�I�Q�<R{o�	�l �U�)p�-l��?bj�����S���?Q\չώ?<0~�