��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P(�7w�}��H+��~ N��8L"�!��ў+���k��`�"f���y}�֐xvT�M���&��%��F�ً4B��M����S`�j~q㞝����_�&������:�|Xӫ��4�;�.P���h"��k��Ԩ����#z�l��/�=.�",hdJ��-[��&�4g#�Xv����ҁ�B���;�s�����I���w!���3��� \��m�#\��Ss�u�AA���%]𜸘quo5�lqy���&�R%$�<��#|�m����a��*�5��c��@�_)pь�	}2Q7����h�ʪF�26w���$$NBn
u����t�i��z��R�:�n(楜jF��4YahO2�֬�G��)��Li�m��IH�j�ft�[C�V���Vv�����E�5�6���w�fw9�T�1�~2}���+ ����ٹ��9�RMR	?tԈ:U� �,�K���kh_�L�Fq2��lJ{��
syEʂk��E^��C_�F�M�rg�A�3ڰR�{@��'R%�0�tb�T�>�7Qt4��Ǖ*��5�͑ �k|,�& ���(� �AK��V�QX:�0}�]�1�s����4Jt2���*g�������Vƻc2D��*�I��!�R�q6;O��U�-�9[jwkO���O��&�/�ks�-\u�v\��%V������)���d܊�6QS ���[�'F)f1�<y��n��7�����7���e�$��O�$�̮��4�|�~��1Î���C�����A��"�����G�Jf1�[U�'?PYZ���B�G˓����	��-���i�
�ە�I޳��7�}�x-��K�*��40�h �2��0���P@Ⱀ�Wj�p%@�S��\�`[CLm`S�u�Ǌ�Vc� �5e([%���,$ߣ;	�0w��G�f�U�- ����|�c��{x��{Ƒ�������?v����F�>A�tG��0ߠM�LER�z5"�嘄�|,�j�m�8���¼�F;�UN������������ D��+��/��s� �m�d��<��&���[ nצ�+�1� ́3}�:���\I��QK�K+f�ö�: \�^Γ���j���G?oF�V��%{���JHbn�̿^"�wI��04th>��#�&gCզ)�6��)6a�䂭S���a����+6��'����(�C��g��Z��Ɍad����Y���Y��߾�>����e�-O��a_�i1"�`��:�.��T��D�U�s�,����#h�t��E	GP�g�y�;[dpu�K��P�n�����U��6[2�<�-8�3c�#I��1+��&����Y'�L\��6^� C���J��6Q���f萩5ͽ�D������~-�q�ƾ�j�=�S��w�6<�`�YQ�vM�,A/
�k���?�g@h��[��7���'�{a[�#���F��i��2�Z`U7{�/")SA�J1<�Y�%�_gR���;����o����)��G�#ƛ=q	��slS���R��/��TQ�.��:y:0?�iez`m�g���-!�� d����c�ț�����8	��j,���>3��8;i����4g�[����a"��M/���UX��uҩ�5z.�_m��]E[�]��Ka�&@o�3�	0�#2�˗�N뫦]��\����V�ۋ�_|�F)/��ך	���R�Tbp1G�+�]v��o²���l�?�4�,��� ��C�=R��o�=OJ����/⏬�^N��(�6��T�b�R�FWl2�v�9���L��ȋ���!v#��l�JN,}ev�j�.�17N���1���HS-ELzyVG�*F#88hh}�B��+��e����R�~�#ĵ�s��O.{���-��\����P����@��Xsj~�	��5�/\���Y�g��ؿر�������6���@��q��ޟuh[ľ�K��;�����\%[B��#ɀ�
?SN/<��
������8s��.�V^'ӄ�n���tevX�I�(p��رՓ�״�'Ҷ��8>��$��1�G%��@FݺJQk�� "V'$��['V��<��jL�����"d2�P�{�7����--o��i�1��Ǹā��O��2�Q�=�e��4���f��J���+F��;S��e������;�l]�*���\;��K{�UA0� �"�䷁2K�O��+��W�Mw��TqW�l��X!�$����e�ό���fg�|w±��o�<�9�+��5�>P1LI�����؈�V��QQR�'�{�8πה������������(����� 9y���,�tqύ�$!��<0)L����U�C�M��3p�lxB8�["���;a�8%s�x (�ǢIG����`�.���w]k���bT���Ubw�!��\�~ec�@!r?'N8�Wo��]�sW����Y]iP�zOW|Xaq�:�S�K=T�_�آ3��}��n�Jn�V,�-h���X�����h5�0V0�a��9��հ���ōb2ĥk;n�֕&p�p�ս�y���u$bp	8Z��O��K��C�?��>˄����.箨��KxuM[����� ��K������Nm5��t�HS�sd�Tm�N�rG���ޣ�E�ڶ"�%����5���.Γ���� ]�I�Hbᅟ5g a�h+��d�j_i���i�"h��U ���Sc����jX�)�-������Ԯ�P�a��]eԗt�X���i!���o�Y�I�E��ϪJɰXr7�u+�F�����l��$1�<D2�+2'ЫcT�>��L
a�v��w92�ʹj������;���XM&m�0�e���G1X���<���d��'�sl��,' \1�1���ft)�j��f|/�.��sc:u�@'���6�����}�g\���ͭ����H��{@��Uw
��uS�>~�&6޽���Hh�	����>(�w
�8)�yX=8,����!�)��7B�Հ��,՞�����@�a��à��ƶNQ��va-�Ez��������߽��MQ����HJ�G��V��9��"B@��^�gT����loG�S�`8�{��g�b�\Lb�z;p^��f�����U���\Ǵ^�k��7~
���أ��I�w����MDT3�嗾E�\u:��뗑�IA>�E#a�u��7��&����d��Ti����B'1�]�ge��F��H6�ꖩP��1�J����𲲗9w�w�}`�����@4Spj�]=\5
�*u�~��f�ܨ������T�	��;t����t���HûF��%D�,4��}NZZ#m�<�.?q���N��ݧ"3ߩ�g����4�@.+~����#5h��z���^�nΜ�@�4� F�%NجY>�ps�LWA���]�ye�p��'� �����R��A��W`���#M��	�,65```�=�䍖���[�X-n�$;JF��{�{э��mU�,ߖya��f��,�������5���#���1�Z�5�WUR�}ky�O���F0�(&HJ�?�8�(G��m�`����g>��\��Z���ܟ#n{����~�)2�(t�:��*a�`���54,Z� WYlX㡹�!��4�m?=�Bݕ[�Z�"�\��W�!�[���~Mm�Z.I%/���5���>��W���Ȓl�H��)O)�!�%�LM.2l�Z������'�n��"Pģ�!{5X̲H��hf��<%��3����B� �6:�%�nE�<�vdn���QR"T�߲�X��&�s�¿ջ ����j�@Ҋ��O"��ݨ���]��7B9d;7�����:%�k���ľ�p�(�{e��E�����y�	=T�e�A�2�aњn�jS�R������fv[���7���!�u�ٽ�?����5�!��k���Ik%�"��:[���%�IW�TJj�e��-pE�F�� ��F��!րP�v̷$ݳl���Ly�Ԩ�I |����!�`���"g�vĭ��@Z�t������j2p���������˅�u�9Q��:R�00�bŏ�D���T�KU[�����+�ӛ"�ѡ������1����v��bW��"��Q3�%\�rW�y~�ǉ�e@f����Q�=8,￧ ��7�t��p�f(5��h�1�)B�:/�EaP$�����]��aQ�]5YF܉oqę$��aZ'��x���=IE��
�*S�_S���u�Y���v�DO�M��>�vݣLy�놓ٴ����R�x�d�֭�mf{=����o��2�?�"_f*���X�X=�xp׎�x�H�G~[������h@�8��R�\= qp�\ i^���Dǣ�zXm�һ�ɕ��E�0�>7�u#9��(c.<C��W?D�E� k���t�OBH��z�*a�݈�b���V@3��g�K�x���'x֛���-5��[l@�xk�{�,���eD�<G(�ª�;!|��
���<��>s^ɀW�߬s��	�����2in� ���|�����{P��Uȝ��5�����v{!vپЇ��|�Vܜ!��Ş��Lod�%X(�y,
�0s��[���kD&}g��T�xט��e��j;S^�~�5��7h
v&�ϵ�5�E�'n�|�6�X�-�U��B�<9/����4��%�
�gL���P8��.�~ְ��jɩgƛo�i��P���g o��n,���
�עf��5���X��%'�7�ҧ������|n>X�����r�"^a�t%��)}ta���y����4�b��RTR�ay&h��Wrf��Ϥdz�V~��5����5�Kvle�B�Qn��P0O��߳��ڔ`�p�V�M/L~�U��LX��Bq�����QtJ0��ɿ�PYZr�eqD��1�\׺Ǟ���(�a{�)�OSM*��?�[ k���JD
)K��U6uzP�t��
Y�zhٵ�r˻GY��V�,]�;����͉R�2='@۝&?���G��熮�}�+B�i��4��&T|��Cq�r�m�!uM<I	��q�Í-�� �{��3j�E�e{�s��4B��Ўn4sk�zW�6^�tj�y���O�4�s���(��N�J����>����SWD7�!��}�h����mP�?y�kX������)6eo5F�n�"��P}]c�Zg�<��lO<f�;�&�|N�e�HN y|K�䐕��<W�y��ގ
�<��q ��
ds���|�bB��]J�X�Bs)�L�?с���Z5��	 "l�� ���)L��f
=Y��gj����t���ΦWE���!�n(���uH3��m�����U�{��CU)���JH`�9-S@�
��͠���Y�I�l0h�C�"#���������ꤸ�l�����;Ǐ��2�8�{��Y�|:����p2�I� j7��~��G������>I�ݎI��ݵ��hܜ�Q�̶=�;�;��=��-���%�=���!v�#�d�""̜��`T?A��d���T���;6�pd�(1�	�S�8@?�xi���S�p�V�*舶�JW�{��d��,�ZLw�wW�=�T�hə{� 2_���O���r��`��
�#��;4i��UF�"{G��-� ��p�閶��|�M|}��M����9��b�cŸc4}8���4�Z�<AZ�X?:C>�E�O�1���~+���n*�qQ�,g���S�V
�Wҕ�K�+��ǉe�L�/�J"k�ux	+D��-���Ԭ|PX���<�l�cX�=P(�#k�G��_��y.����s琹i빛Śc��h�v�{���^]��K:��e��xX;qp��::���&��1�u;�FW�Ͽ7磙�I/ӝ����K �O:�}�����[=Dָ`�O�7ܬHm�)�W���w������~��v��s،E�֢�z�9G�n"�y�9�imR����@
�WY٬���
=fC�9 �a=�>��S�A�B�}@"q�W���q��Ƃ�����5X�O��6Zw�`����~�~�Tf�o<��B/��b�[-ȳO���[�y�UR��������a�!8�vK�cvB�sXU�k&}a�@���&Wr�(:s5%w�h�1��g�g��~�J�+�Ҕ��J�O�� �=q�C5 2���@��ǔ����ABV�pTi+����;J�&��忺(�j��V��}92=��p�A���A���,��G�>����o�^[͢�ˍ�F���#�ZB�jp)a��p�T�����O���GMF�8�Ǡ�I������]?�F��#��⊡���PO&G?ΟF�i�c�y*QrIC?6`$nO�eMp��h;~�p!q��ИV�X�g�R"Y�ȓ��巯Z3PGݴ�Ì�I���N¾�[�1�^J�57O��+�s�UX[��ukC��g���܉���(������[���|���(��T>i�_�gP?�k�1��#�:�.4��b�� ��(�_c~:��\/����JL��/��/E�UC����t88͎s8�m���f@a�ЪR�`pDS�_�b f-�9���w逓1�T
m�ǔ����F��Ff��$��E;^D�1�E�FX�a�;�2M���mq�i�x��:���f5�6�&̊̉~cZ��o���X�Uh��Qΰs�].c���ғ��D�>�"�����2�5�2ÚP�`/�m�ռӔ��7��5$�*�wm��"���N�1��1��<żUг�%&�8I2�f�Xu�h��C�;�G��c8n�z�@�1e����;���A���GO����Oβ
-��FvFˑ��lA�`���}v�C��(mUؒ�Z��f�m��f�r#�����CrWiv�-�.�-W�Ǘ"q�xa�뀸��l��N;������>̎�?�˾�y-��C��d`N;LB����;/�g�o�->��m��Y�=��L�q}�4�R���|v*��ơ 3Z,�(-ϞY�o�ht?��bQ�;��j��Td)N��*(! ٭m3�,��Kۣ�+�j�p�O�X����An��p]�Դc�k�s���J��M%�f���``w����y����ʞ�ʠ�I�F�o#E��K0p�?��(Y6�Yl��*x	61[�Kz�Ě����uY6!�s%�?w�oKJx%��G,���_�ԑ��w�3�H�4L�Z^�U�E6�>q~9n��3��u�9_�ΰR]T452���0�&t��P9��#vM�����j����r(V=;�s�4p�O�Q$�Z6�Eb���m ��O�[��d-��m˔4%�M�7|;C�.�5 ��Д�K:"��:�ۉ�,�(N�M�7���I����z��|gPlz�X��{�y?*0+*�]� E�����oG�����-X���&	��DŢ�qg"y����~@]���������/�pӦ��dx�i�`.�(k�(绮�h�<mj�YMr��Ds���u�C�Cvg$P���K�I�DUq�Ԯk�īh�I� ǣ33r˺���;�����${���8�Y�������� I�'	�Μ�r��/���&�������}E@@�����g�qj�%
�#�q��@v��%�/p�5�P��lu��ꘞ�7�D������{����Vz�"Z��n�[O��"qn���+�%ʆa��Q\j����G
�`�20|5_�f�6ל��8��t s��,p����ZA����j�%+N�Ԟ�Xʢ������
�a:��iE��)�P!����g��Η��섕��ɞ�E�ק5����H���5��ݶ�}Q��T� '��LRbx�,�\����>�PT�!9tA�>���
}�J}���O6��"�Rz$߲$���̄��IP(��d|.{p����o���~���F%��K/��F#�f2�h`�����յ��3;7�B0gau>?��17nSm��y�O�ui"_���yTfЬU��>�s�)�-��kx�]u>�K��H|k\i6jx����ᇤn>震�Z�U�SƁ.攫l�'�OJ�QfV�OT�����/�;���z�K?L���,���PH��o%�4r֘�-�8w�����>�SjiI_n�룄ՠ��x}A F����P�!����� ���J���R:�����Y�]��-OE����gҝ�"�G�\2�c ӻ�,Zf�w	7P1J��gs�ģ�T����?�ߌFNt�Kl�KfbD�����L7��b�ud����=�7c���bW�9�(:jLDV���3ԋy��(�FS��!�O�ٳ/h�4>�Y�-���;�]�37�ެ7|Ηwzh{�����E����T�τ����U�f�]W�oƣ�����'%/����r8%s�3�6��d�h�d&~�iՙA�h6)�P55.�ј[�|�m�
̒��(��~����*������$�kM�m�}���5��ܬ����%4�/�\������LcS^�b����/C�c�ߊ�|��`�M�����D��2��>2GY�j0��V�S�"���f`�
|!n;��SL�[��f���G�ל����3�}=X菛�Z݌�_�R����帀G��^�٢��r7�$���*۱;�o���5���<f;�l�"��T�o|�F�v*E����`C�n$ΠuQl; fȹ��]ۆzb�C���`k��{ܙs��G�p�)A\�_� >�GH�I�,�y+��T��9ʴ:�)D_���#�x�`t���g�j*::��34V6oZ�Bg�C�=������x������R�A��x����ڭF����Z��:������`CK�ii8�+�	"3q,�w:*[�-h�]&,C8}���ǻ�	��'ٸ;�wV�eU�����pw_��� ^H�d_ϊ҉�9�$�I;��D+��+?�]Vr_r� �i�ma�i*s�J�s����0�S<ո��{�C�A��$�n}~1
��g��Fx:��� 
7Ŭ fr��7�6n�.�Ե�JwX�O��K�����#㏫�Q��;�/f34��QnNUി��Ͱ|�邜X�n��QQ��fcT��gߙhi$��r����o��U��2d��lXC̽�x}��π�����^ �<6�ʞ!V?���e��2�w��cE@�y�BIi�G�pɮz����؟1�z�P�Ȯ�z��k���gE��ca��1�-��Y�?ס�R�L&hzj������p@U�劝D�r��1����Ȧ�]7��#�Ҷ��~�;~*
k=q}0�ײ	�¬��s��hU�{���ϊ�:*���vЎ=I���^�
:��M��S�AE4�$a��k�hl�馒����93K!��������f��RK>�3�8��=���Z�3Y�:_TUw"DԭIc�),�Y�4)�VQM��u�.�K���~�*�yV]���A]�28*D�h���|���*��͏�p2j�$2��G��h�I}�{œu}��q�A~�P���[�Թ����i?�h?�@���s뭾I_\��߲�����-��i��KA��L���ű� ��^�)���j�b�w�!<�>�'��2(9$�2�v��Rz�@��"������E#�t��F�<Q:\��XGs�1�g�^,;��J
m�X]�*;QW8���ͬ}�ekHv���Ě�Nn)���U�	<�*���
��R��B1c�j��{��,���"�_w�U�k��2�F5�J�N|*f��f�3�����,K!��M�f�j�$?Tf�<��X�?!���+�5;�GD�h\���B�����VnU_r<g��E���Y�#r[j]��8nw^:�.���PFq�)�D�5����!HP��§^U�D��D�� ؕ.��xAҿ���xA1��#��^��1�����R�H��&�J�T}�����ڽs-.v,P)�ST]#}��v��)�w���zZ���㬞�Lo&.��N��J_xB�� �诏iཱུ/�vEK�a�}o�W	/��ц�yE�۠왮 J*������f�?r��,4u=�9��z��4��.l�,,<c�LQ���:k�/��/ɚ��?�D�2eY�����?e`�ch���Ff��%�(ͪG̠�	C����F���V��Ea��c�⪕iO��,�b�"��]��,�����3�v��_ ��a�"�Z���]6b�=��}+��`��i�*�����";��S}��$����k��_�c��Q��Q`�k���ts��/�)��(����N�@ٚJŸNyP9�b'���&�m�ΐ��wv9<#�Æ:m�?��S��Ȩ�<ҥ�V�?���z��J�0��S{��Ȩ�
��
	(s���8P�j�`����k�J+��؄
�ԨO��CZ�Z�yJ��AU��4��_�^�{64��J6� c]�!���~�UK�a��8��6�>go��df,�3���Q�E����l�4�u�:���a��QA�}W\���RϷ?	Έ�2QrgO����K�Jq>S��
�ͱ�YG��(k�����^�����~ޤ��j����w�!b�r��a���j�~����qT�5��� L����O�5#D�f�,D+�GGG�o U����,eV��IZ�������P��w7H���=h\�_�)��)��a����򱬖6��?w�]�K�0uV<�-�Z/�8��1�[��2�
�XWVb�g<]i;:�M�1A���u�9.����/䗜4�wI�2��R��n���䵳�E�P󽧢���I���w���"z��Di �-ŔJҊ�e|�@?���������.�#c�!�x�7�+�?:�T��o�
o{C$Ƭ$o�f��ϭ�����j����z�;�7Y�L-��Ɵ~'bٿ<�t���o5}��31&�Q��w�w���?���c���t2g}?�\�g���2��U���X;'XҎ��C�
r{��0	O8��JG#h�nim4����y�;��Ep�����@�Y�<~�!�7a@ޛ�* -u�U��οH���s��>���Fu�`�p�8� �5�H�&�I��2	 �*��wPզ��ec�ǀ`}�X����<�06G�kd�%Z�<��N�5�0�����,8*�B�,O/Ӧ�d���?�[\��\NXG�&��� (0A�;<��%e8�)$��jD+�[�f�D�]u��j~C0=�7bW�������7��j�,b��XZ���g�H���)�M��['l9eGV&KJ���ͽ?p�i�9]9��l�c�~9��*)i�E�ݖbg�s�`�UW�3��Ut��t����_�Y�E�}A���������ʇ���lRzW#�W]��cܶ��E��}E6RE�4�	��)��v�\#<��2��~�F����b�y.�+fV��r�F�S�� 9�������a:aX��(460ݧRc#����X>t�@���&d����"���,�?�#�k�|)���
���N�TP(?�r�O���
�x�G�G��N���fG�����Զ2-r����;��������Y����a209S�vN 9!1�� T?k��x���\ӳc�ڔe�z�S2���A�c�/�7<�S�bb�Օ�3+���A�4�n��(7�H�ݖݕ�.ԧB�����1r	G/�6�F�̹j�\X�:��0�њcC�����4���tڋCN�돷�\t�F��/~'W�եZg&ֺva&.�P���~2�5�,���\�Μ\%~9E�ƀFZk��4*�7��N�jjV�h�n���Ld1WB���Š�=	}��No*[��V����Y	T53�u����#��$����L׎.w&)��0�v�g��)5�:?VA^u��[�Q(�α�����SJZ��(�--�����?=���4�@c'_s����r�Q����##�hi�1TPe��R��W*��ݾ�Y�h.NL"������r�j��fd��|�]f�F����H��J
S5h-�H�����2�j��%��?Ds�Ն����!K�]�G�Yl�{�A��fݪ�xleE�-������o����C��,!��3Z��A���0�/ߤj�N���Gq�h����i�p�$I�._�(��
̙
҈?�e���U��Z�]#�)�X������i]�=?�j��fJ��\щBF��&S��
j-y�$z�C�H��}+A49��ߔ��m�m�K�+��d'W��+�Z'�2f��lZ���߯��S˰���.�)I�'��Y��:��։=�T��� ��T>z�q&�Y�,ڌ�� 3��A'�tu#�0Ѧ�`���D�2q Y��⌕�i�����=�9x��}!�	m�j��IU�K�
:��� zf!J�P���т&M��9�||fn(�{��W�����"N#�ɖ�!�/��99ٮH4E���<����x�Ky=�&3|n�E�/��� ��#>�-���T/�+g�CdI~��3��q���6>4��2��8�W�@�뤖�+n��\�4pu^{s������TP�{?���P���~���� B��qƺJ�3mցIgv�L�����5J:�ÜL�Hq��z�R.��C2M�cS)1�t#��aNr�uq�������ȑx:�;u���Z����p��%�]��kΜ��� �P�5Pf؉!�3��>�� � U��Y}g�to�%�D�oy���jtW6��,�����>�]e��!���h�;3�q�io�rB�P�-��t�3 ��2Cz���k����Ј����a�],OgVG�E��tl�ӄ(׺Xj'޿��=2TQmB�u1bm���&��<)�ב0�e�ɟz�a�����u�g�'J�O�#�'`��!����q_]�V�&<rH�:�a�����HP�R���D��ueV;D�#�ػq�"�祜$�_4Z�0{�Rt��kk�5�Ӗ�&q��z(�KYp� �3�Ê(�I��7��m���]�6��x�Edq%*��?#G��A�pF҆r��y��M������A7d�,������}�t�Z��q�%��o��(����jA)�t^*��2�tHm�*��6�~�(e9�6���'����n)?��U�O��ꎷ ^���:�yi�o���^���~�I���Ǟ��fW�\�Ȗ�4!
�����)�=�F�)G��[������=�=�	�5�/��]�w�:O�:�����-���Ej�;v�GL��.H����>�TE����F��7����~%`i��>;���6�IO2�$8��Q3��v?$��(�`�x��ā��n�Q��/��oƚ��@���ydgк�+�9��r	��Uh��I��1',Pq6k�j�GN�B��"����n$��l�>�yN�LoF��e�%:����r΅�6��J2R��_t0��f79�-A8_r��A��1�.���!��̼��T�zh�c��S9X���K��<��0ٞ 2���p{�$����8S�dD74������M���~�L��֜/@�'�z>�N����kRs ݡ��w�M�R �"�'�UU��RD[����e/l+)�������UW��<�L��u�t��Z�
� ċ��C��*|�D���b���0_�_$��>,���H���_�8�$�v8��m؄>kr��7�4%����mmR,�,�=�ځ�D���6T�!�{)�4,2��$���I���DZgO���ܡ��8�h&���$1��<�9J�`c-�h�k�F��iOxM��	�A=�Õ�LG����Ϳ-NX�,K�w#�:ً��v:���eh��χ�r�:�[)z�̱��t�ŨRBG�wG�6��4��׸��^�.9g����nl�ý� 6ȶV�v�:�qB�|�x��+���[U�&P<`���΋�G�v��l6��'�X��PT[���X�K �tV&�*#�#Gå����t��h	�g1�=lE����`m{DJ"G�+���Ņ~�6��OZD�8KGI[�:ʥ ��`����YS�7�$�"�#�*_e�ƚ�"Z�dp�᲻s-)n��Xz��~A�/�7�����uB�@�yȇSG�\�����=�k�����瓡uw���^�,W�'��m����9ǲ3򔝮9��r�}	y�����s�4�o��)*oٰ'�U�[�SczV��SȀ�]�B��ߑ|3����ܵRZd[<%����a�̶��]?>@��z���0�4��M�ܒZ�����NC�)���gV���J�p�6���{���>�'z��.� �7��&���j�^����:W	��!�)G2��X"��o,y��9��¢�H�&g���;3\F��&���`K�M|�"
��ղ?*s�#��g�������-�,¢GW�ѩ a��V1�2������b����p�k�0�-xj�<X���ݮ�Ñ�o?9rL�9�a!U�6O�8��SїX��D�e���~�Y6m�� r5�}u>�
����{;@p���e<���Cf߈��W� ��u�M;���olץ��6%ң�e{������Z�O[V&X����6��p�h�%��w��`5%���[Y���fӃؚZ4e	�F���Ղ?b����*&�K͉�\rFF-R��<H.
�{��C�C��l����e�K!ID`��M/��E&ag�Lm�<���nZ����8��i؈c��)�_H6
CKF�7i�F��d�9��EP#��R��-�5�����z`)��T��-R�'@a���_��}���J��=M}{��ۄ��w�K���,;,X�&w�_R��e�)��Cp��`�D�'��][`QE��D���y_BmD�0�s2H��a�X���^}�wh�(	G�)Y����a���d��3]T���Z_4��WO7�xr���=�����ĳ�m[��Ff^�r�.��՝��F��/�{S��qA����`�*�a��Ec]�d�_�|�Qa />N�����9}�>婹�=/ӓJ�Y��V��H&��˪7`�Ɯ���9���|�5��
�_�dtܗt����֚A���������A9�l0@���lA1�U�;*���njX�����d�.�:_�Pi:���˭>hhP�BC(��0kPgh�<���"B���� =iv�5�����
�p�&eU&E����R�^fv�>p�Di^?��Ed�8��C�:���q��PM��B�n&8����UO�U�&��zq.��z;3�2l����&&�ĶY^�	Ա�����W��������t/�M�$=}2�e���Y,<k�|~b�$[�.0�Egd�8|.C؉��i��Ao��v�k�mA���9	����r,�ë3b�#��nC7!ޡ�}h�|��TB���j�x"���1O1q�8�����v�8�\(�]��4v����"�Ϯ�����A�٤�� ��Wۛo�Z��Up����-���ؑ�)��ZC8C�U1�j�>��chz�EN�B���5��](�a��Pa�0�T��1�y"�V�qQ�Ӎl^ 9%=#�4��<O�� �<�C}̮�!��!�#^sC4�n�k@��Y噬����� �%�<;�_M7y�^X?i:C���Cz�ni@V���+������B}v����W]��c������cMU���[Y7�PhԺK!~��.�X�+ҭ�p�l���j�U�dh𤭬�C^�����R9���r�n�w<q���P�!?S��W���ʴPJ�A����`�F�׿)��Þf�o�9����B!\gD%{���@W/Q���\�ǖ������7�˝��U>gKc��Qp06�ղ�;�'W����j�(�>����_fw���}��>xp����t������?  ÙI�������H��BL���P}�s��Ne5�'�{��s�^����$L�����f��\ay�V��T�%3uV�R&Y�fa�/(��ML<_���KmT���))��78Q�������Z��<�����K:���k:^�+�`��^nQ��$:����2��k:�5��5�Nq��2�d�E&�u�6��M�j*)��d{kI���zQ;X{`�eB�w���ʣ3?�> ^�g9��d�G)�/�4��*�BF�#�>z�|�
��u�B��Ws,��8Gnnm�9U��&N��[W2:+،�����@."�>��0���8�sR@�'�R�蠰�|�C��������z�z̫d��M(i�8d�tzGDO�& L���$�3�-�z�Ow$�Z��Z��,a��$b����({Y�b���<!� ^�'�ֱ�2������%	�#j5l��A��A�}�3iC7���u,��*�\���[��F�w:���%8 z#���2c`cn�	��^"k�p��݆9��_*�*ws�<2-��t^PH�� �%_�'"*����WJgT	�'̄�/%́@�h�U�Ę6fA���I�(x@C����y�x��N?	�8��Z��ps:���.�B���K�����n��ꜹ���S�rO!6!5��C�`�%ۨlL5R�EYrS�s>�o0J{����(� ��n��0�]MMŨ)�2MXM���a���Z�z�e���1����d�]���k�q��1!���$gsB���jD,���\�b&J��gǜǮ��/yR�o�~r'Q�t��]ަm������`<:����
�8P2�`��h�u_�,��!(,j�%�M2�b ~AF��k_Zc�L�m���	X�ۖ��}�OtIgǓ��/�'5W�Z�m��F�E��"�K����YJ�����U}5f+������Й� ����+�ns��B�E*z��Y4��F�UE�́(�=N�ê�U�*`�' Mb��ffgP[�@�ez�S1�I���;v\�n5���>��B��^X��-ӧ(c,�v�۠H��Q-*彡<I<cq_؝�ns�&!Q%+<���!7��\-����A|�l!��C�W\r�b/��E��hH�	�*v�1�$�@T�҇܆u �b���ROpBA:��(J!��À@�c��+�q��ٱɉ�SF!��"jR��}���k�߰���BF�)��St���N�@"篲����1F���s>e�������Ud´b�o9�K��N�(ɺ�grkC����Er�F���1��k&}��#��ي�{C$�wq��¼t<g�t�:#�>�H~���!�o񲔊{��WX�\(�Zu1w������t�,8�!z}�x�:���͕�!*�	���dsN�ej&��#�l��1lD�!E�8\�#k��R��%�)D2r��t'zj�#��K�b����85U�R��	�bBi4y$������=\p�
��唙�f�T���5��`��K�`�eH>u�,El�D�m'6@��9$���H��彠�S3Z���h���oYjb퇡X7f�U����q�����Q0G��L�+�T��ώ�8�Q�bd�gU[�U�9�sW�{*��H=atĬ"�p8qWq.�n�gSq���~l�ec&�取�Zl��v�]²JU�f��!���u/��De��ԁ��H�)+�輲�Le੏���@�wZ46n�
I���\3��qL�|���V�a�/ȃ�|�!Z;,'=�s�H��Y<Se�jE��^�w��q��8j����v���ڱl������F�&�[!��^An��'������ܳ%�u�w���@ ��3M��Cn^H�֊��
��,�Q�b��l=�&��=�9��n�%,Q�w���^�uVm?��b���7��3wR�>c�Ƈ�`��~�-8%�m�5P���D�V+�i8m����ޙ�yжN�
#�ĸ�-����'�Ts����)�>B���l֝��z��ا3����}�7"���D��Nr͎D����)��3�K7�ܧVNY=�/V$�YZ��߄FNƪ6\�c�� �-�/J�Cs����8�G3�SQ��0��5�z�
?;c�X	ye(�Ϯ�g�AS�yPh�RZ�n�MJ��a���rէ^������'��U�-�@�]}++˴��f^�켍@�ig$�N����E�x%v�j}i�@l0���u3Ģ����7$���T���G�O�<�|S�)g���:�f5�Ix'�\/��u�#3���=��I��,��yA�	UOE��{AF���
`g`���b���b��mz	��mw���N���Ɲ��k�W0�T���\�]K���e�&�?	>�Kha�ju$�;;y
Bؽ3Wo�R]D}�
�.�j�r��OT�B�=�UK	��[�Y��'R%W�<�����UH�+c	�kq�0�����~��(���۪ݸh��ۮ��.��A���~Tg���R�U�8��b�Z�ﬧpdt�4�7���+�c[��=����GQ&�  �F>�ʲ��Į�@T�cI�O�d��(�ȬT�4b1M\n,��?I_/���pF�ݲI���f[]$�F7�0�2�aZ�W����v�Ȏ(�+aI��%���~�MNLu����� c�
��EVd�ױ�)��ĀQ*�� 
(y\+�̯�����2[��p�2\�$��xuK��.�!5��,��+O��u�p�:���/��9��ƨ�_{�:P]C䛖M��lo�+���գBť����Dr��X���ʽblO"��zk3����ɮ"{կ�r}�J=]Ɨ̮H�Lų�41� ��e���
`�֊��y�8�=QB�!�0������,��B3ZJJ�<�g
Lo-}�ڸ�cqOΚˌ�8@���e�Uπ�^<�"r��b>c���N�p&�?�ͩ��ў8��}@	.*P�A�]�WI�o���P7�'��߿Y!��H7������&�d��^҃>H=�h=u�������>0��� �1`��|j�E҆ǬDBE%Q!�l��$���f����um�n��>Gx�b�>�[+��^���
��ۏ�3���Z�E��_c]-;)���G�����Ӊ�:��z8⼴�Ie��=�_#,[��T��?�	��TT�k{6{��K��axܚ�.�V�}׻�y<�zY��;���裴�7`�'ټ�40FB��_(sS?D
h��bp��i�F�ao�b��r��l��H��:�:��z7mgs��W�� 9#�9΁67u5A5��(9�E����D��j|C�:,_�h��V���t8زO���GL|�μ�b���p ���!βȵ1����-$k�u�)�/���D�c(�wp�og�����Y6�)8���ӷ���2�(1"�x�o����2-Z��K�ĵ���p�W�Y�'����I��}�e�����x����l�)8�L�"�>�f���D��<�}컔)a��8��>gTJ5Aަ���z���&y3�=�.q�� �~��J��WÇ�����#��h��9�Bj:�B��XW�Y�1xȾ6�w
��%���!�x�@�((�[���4{�2)��R��A����Kjh���G@��)����JZgMlQ��!������g���Jfx#�.��[�6�я���~m��Z!B>?=��7�(v*��[�%��J<��A�6�,^s��9�sja�q�̕0t�q�w���V��6�(���w�Y@/��+�3'�:|�)�����{bqj��%x��Dt��QBF���?B�����Cf����*2���~v��*~.���z�4R�\�M��hDd��݆5��Q�q��:EM��`oMJI&��KL�z�NN#�}����.�vb�~*��4��YM�����m%|��
5��Ht���2Y��,�>lV��Spe��/���K50ک���?���M��m�y&ct ,��ETv>/�ِ���U~��(�A]��]�G����y}�^���������DvS��B
�$�Π�=��)�̃�7���K͊�Kd�:��ӇO)��&{c�o�^�f��۩Ffn��>�&R�2Qn�K|�a����0*�A�����Q�g>�Y
h��m�y �V-�g��ꯆ��5��;*�����43X8)^�	P�f���6җ"�֐UR[�W�\�V����w�:Swf�?�9A������(vp5"B���9��,;��r�c�2uNN�a$�~��^��T}�4?�5��^�
�݉5U��C2�\#W�M�U�ʮUSk���a��N<+7��;�|̅ok�*�� ����}�~esT����W��PAiHWi�S����߽�?F�&�?i����8�5�ӽ���Q�������*�\�MaG��As1�e��3j���j���� N�LC��d�lDh5!��������)�M�aYF��٤>ӷ;/΅ Ϲօ�-���e��$d�T�aF��&" ��I��'�Æ-�TM��s/�1�'�M�T׽{$1��}�z��HI�1�?�&JC��Ϝ)�Ì[-W*z�y-(=.�8<��J@W|.K�8�i]Ja�u*Fׅl�䙰�7t4���tf��W�i6I�(�-	� ���|�g޷�9�v��h99�C����n^$���*t��]*V�2D?/���B������eĂ�
M� [H~�x5�f��i�lF��v��+[.�u�l��˚�@�v.�W�C�Tp(�K�R��M����CWHm@ ��3z	@��g��a���Y��¯�?�f`���>1ҬM(W�gV���ƵX3D�@!:{�ԼuX��+D/)Z�9C�H;�����
�Jp�B8�e�<.N��څ����Jߗ�Z�I���+��	J����;�ͩB�z���r$��a�ځ��˶Ï�W��u��r�ϔ�ۢ zj���� a%b�����H�r����׫r0J���g5�D�yzO<��.�����:��җ��W�������^�T$Dy�.GoD�G�fA���킾w;���u��
]�cӞ߷��3�t��3  �ג<�,'-q���Q������&��o���NEQob|�%�͵�q���\���	L1����=�dh���b�A���/�y)�
S-.��Ԃ�s�y.��W�=B|���+d՛�]��� �����c�7���n�/$<D�#���C�����(4�Tf�7�}� U�y<�y4؞�3h�vg�;��x���HpLpG70�~iL��|bP9@8O��&�� ��KGr|K\�ˢ�~P�T��w4o�l�d�%��}֤���k3/y��g�WǄ4��r|
�q�j���j�}��� '�1�CxH��S����"�pl8�[V���TFo �F6#�!�h%�^��"����>�y�>�7%�ƅ������
��dn��q��C%.Y6�f�L$&�|O[�ꋴW��  /Ra�m�Bzi�����#��c+K����Ӎ��A����I�[6�|p�YQI��8dD��0̾�5�Թ���[,��\V��P�%_�)�&}�Bإ[m0�K撪��X_vig�a<��<��vm7�n��Z�cޜA8T䊂�N����f\��\���=��/S�X�������j����[y!u1ܷ����M�<{�H�h�zW��aȵI�{�h���w���㓢H��qA��ib8�J���PVލ�yqrF!�w.�1B�e}����±,�}��z����6v�#�؄X���������P�����<k�Q�����װ�w�4���6�2/�*�j��%K��[;*=.�y�xu�	A���vl���^p �� ~*鞊�tD�����Hmס���zr�rޙ�����H�����.�0��@������S�l-�z:N}�`i��(t)�h7�����{Ċ��d�Ք.AR�.KX�&��e��oNrZ��*D���8��1!�%ߊY��|����ĩ�#Qm�XI�y���� 4��e��m>W�*Y�d��6��f+e},7�k.�\��l��%KNP�ᴱ��x�x;;�#�U��m&ET�!8�Md�j4kk��P�m�b8��;q2y��@��s�!�W&ϖP��` �ָk�ղ��(ǭc	����'��!���"dLS��}�Ѝ� E8Y�ļ�A��D�?S�1�X�����;��\��%=��_���%����9��:T&Z�E:Q��.pZd0&}���m�MZ���+�Ի+Ϛ�$O�s
I��xGN��qǖj�k.�[�i��g1��ٱRΧ�?�|M�6e*d�"	�v�P�d�q��!�<i��j�_3��k����6���~�8�;Y���,<�4^��������Лޖ�g���xj+U:F����mnT%��b��=x.�Ex�P�M��*�$��{a��e}#��g�����=ѱ;�:>D��:��Q���7)�1������.	B�,7�^@v��;�i.:�|�n$�H�ueї�m_����C�1�b��H�6�
h�8�i���iyȝ٤hq��SK�¾�ls�ѭ�mr�R�N���	<߭+HƢ&�m�~i��Sk��P���؎�J	��r�Y�$%�#� Vob���MFX�	�kF�:���l1l�k�S�D^�Ք,D�}z�?/#�o�k���6�C��I7��2j�U����+� &��Z�h8� G�;�CM�]8s�M���k��H������%�$�x����l@a���t�sNHP��g� ��Rq�|ir��f�]�����<�@,v��u��=o3���Ʊ�p{����������v�m	~6��$20����_�\��1���s��1�I���ʏ��F}q�Ѿ>�M����e+�7��v�s���s|E�zEy-�i���^<M�O���ֱ_�m���D��"U{ݝ��zz��΋j��`���g��̆���|�T�zȥcx���~����ζ��?iŀH��
���ҫ�

�FJB����0	tb�o��?R�g$�&?��}�I�J��9���}�5r
�L)'�����2��L���Ƭlf�豂���! �,�dO�!K��1����
� ��(�aFT�k��|�2szn��$�ڞ{��4K��ɴ(Z�N�r��{�t��1zRc���௅�c`1��+�	����Ť�BSoU�W��Xv3�Dh��*�8[s�ԇI��v+`{
p3�Ձ�^�XCfkl�i�,ØQ/ �ݠ��Xq��Ϳ��DV�72+G�;�_ �x�����q$����8��;�J��dPCsC*�j�i���#��Ty�"PW��9����M�ytp	=@�=��²h�vqD�����tYKp��Q��f�0{@þ�#H}�b���7w���]���f$_�a�i��Lm!��6�]�=g���1�םҍXBB��}[��|��V������@�����ay�KJ������E�0ͦ��L|���bʨ��{�*�x�C���í�YcQ�*�����\�KQ`�}�ո�U�8�Ms��r䄬Ko9���"�5<W��[��%�[�L�.K��9����sO����ƶA~_kjj�'�����J}�4Z��+���
>Ł/�[;���]}�s!3��������v�=�I�C7S��Oi"v����i���S<qm���΍��XQ��\*�<���Zƨ)'D��e�t\%m�&�8	��R�!eܒ�{PZ�39yH"aҳ}�@,�0v���b�s��ݴW��~'���g� ^�@���?�2�\+�-tQR� �iJ�z��lI}�������H� MP���.j]-"/r��^�}}v��y��T���($釘��8�U%�
�q+�S�K��yбZ��2��P~0}��f�Ե~O�I�N�\����/l].P���$�њ��!`AC&mp���+�a���?�P�~�8g�	!���49[E���$�#Ǳ��9��2��`'�� s3��Ѽ*EBt�	7s�~s�v��4�-�R8%�Y�G��3.���rw�|`���>��ς�Aj��� �h<Џ�&�.ȝ�T��r:��Z.�N�k&��T������Kg����'���gɕ�B�ً0ւL�xMh_�^KEo����=n/�i���,�͒౽'�m&j��'�3�	 �����0�o\b��d�-1���V��A
��G�؉��B�b��3����L#��Q"��ԀmZ������p�h���tY
�37-��e\eF�B��-]���d�b�0Pv(�l����s��V�236rqmҲ/��s_1r�������W�ru.A�^��Y�;��dh��+�yMl�S/�ӿ��+��}�ݿE�A�XCM��z1�{�s_����-�^� ��]ʹ<h,'
x*x�.��7>5��rTߩ��%M�6��TP�Ū�u�&L�h$�f
��+.v�/�_vKSa�U��ek]��/{&�w�И �����a�m������@��y�p���h��9y2�[[>�%1X��t߅bU�Q�>���������Q�p�&Z9�	S?͇v��jh7P�>������L�v�o��1�����G:q|0�s��g��C/n����l�g&� �����
�x�R`aye�������!j��dz�B,��;+Z0+c#�(�⺩�S������gPл����X�}�"���~�Vʖ�\b����1���0�oҽZ�_73���U��c�1�Ѷ�D9?ҵ����i`(������Ha�	i�t⇳����j���(��6���Ƙ| �y�{N� Sų��;@<C�s���Q����[�^��n���dYQ�D���/[7�[(m�A���v[���� r&������XWź������B'�4tq���D��t�'��-��Pm4)aS�H	��*#��v�p��B�����NW�bޯa˭K�������%�/12`Zb.�L��u�����Ʊ��o�^�F-��O�/P���f�k�r��M�7���"��	�s���x�r�{��#&��?g��'A֩���ɏu&$�tD3#��}�o�E�zE&4����Yi��˴�q���-�I����Ԟ������YD�B�Rcu5/߹�ri��F�ݫ�XY�	$
Ɲ"����,��C�������<hC�yh4^��p� ���n�q��Q>��ώ�V)�F�"V/|\�SjH�x��/�H���s%=��p�wܗ�H��a�|���� �J"���(��%��ya�ݯ�͵M��`�;�U4|V�8�G��Ť���>7@���N	Y��q�>��n	� L䎉������%u�NNsi�b��dV<�d �)��S����Jb8�,&���W!C��~d�w��~�g䘣��˙�K����m��BP9VxC��g���,��z��䯄��#R��"�T�;�*'�MU3����(М��������q�ME�<���+M�g�D�x[ݚ ��?#���Ji���@�� d��]�4~;�Ce@���}�l�k���A��ء.nF`s�*��S�����-%��1	h.���3�`�3i�=�Ŗ)=Sos]W���� "�d�eBS�	�E0�/hs�n=Ht�LUp\�F��<	�ұ��� � Ր<�hUX�X��X	G�$�.d�����%�*kl�ai+���'>mA_��B��ܩ)�BIEI�?Z#X'���I&̰>�!����|���aIU6чSm'i��l{���"̔0���-�����t4p��t�F��̐ԸJ�j�A�^7���$O��WC?W�p�������v���!�}�㎀�c&��E@� ���(#U���9�v���ukʯ�kP9���(&=�?�\�z�5��>�������F%�W���q�k�b�M�P�^��� d�@���?�֠顾��)��� �H(���e"�Ci{Y)�i���))~Is6�ӣ�Ǯ+�^��t�8{Y�e�R�-�䐤�s�]�= o}�57RDw��	h���pxϺB��B�X!�}���-� .��x��e�ӧ���Pn��97V||�,�	���Ao~�47/���BM�i4fL滚r��7�t�آ`������ģ�N����?�n"s���K�i���%�s���Y��N��6���K�o4�:*@ܯ�i����GD=U�g*���	u ��P,cQ�ژ�}�Pfz�����U�2dl��U�$�� ��A��	5�%vBڟ��pxOd2�&ԏ9�͕���
ܫ/�.P�{B4=�-uPO�-��.�;�	����2k_���R�~�U}͐~B{����0�1q5D�t�p�G��ΓU_Bk`��g�������?C�m��bq�_�?Oc�;��>V�d���4~���0��e��*��x�ŽJ����h\����'�ks���L4^��s�Q��P���m�����V�Q'��I��jk�5VJv�rLJa%�nr��˟/G�H��"�-;�o'�O�[�X�Ǵ��7�C��Z4��0T�?!�D����u��"X,6Ƣ}�/J�`A��݀��������F���e"��-tA"ߢs��Rw�Ug_�'����).{�x��Z�2��%v��鮳1��o}eoz�����dli8�>`�x�M����
lb�:a���ӛ�/ml}lt#7_�h&��npP�9H9!I�^5�'��w���w��wT���h���|�˗%���!1һ!���\�Y]U[V� ����Q�31|�6�8n�խ*�P$�-p��o��� � � �X߳��>�e��;�#C \��E�;��q2b+�k#���~��_�C�@����G���g4c��'$��y!�Ȓ�i,�4f����:c���/Џ-�>P��4�/K�u�Ֆ��;�Z�۪-��k;Ɔ��4P����_�fu{b�nh� g���蓵doʆY�Rb�TH�j��ݝ'�X�=��L!���7�1)=>b6�(���U�&m��<*T�Q�p���w��w1�s����3�6/7��D�k�O���t�@�8�\8,F�c��+*��`�)��^�$�XH�>�o6Y���˚������|:&��d���gb�����m�I���ě[�H���?�tz+K�4&L�K?�Aಕ�4���扲�C������c�J�t)�j8l��ȹ���NO��2��.�#\�·�h�p�|�4Z6��`��O)�S�S��DN��z�۩\�V���ҥk�� ��?���� 빊�E��Xv�����چ��k���	�M]���ߨo�'�V;
���P���-H���2���[��y�t��Hv�����]M��ܝ}N����$
 y�=���㶱}�� $��-�>��ZN���g=��5��R���N�b((kS�v#�L���q�Y�2��
�t��t�Tl�R^�7Z>�� B���$%R�r���p|���3P"|�4�^i��O9�TO�Q��K�X9֥!���V��Ʌ�Q��QF������y,ѣ^���i٨�v?3d���� �у]sw�[�J��u.���u��v.�K���d���� _q�S
z�g+�X��(�ZoP'}�Hc�y/��k��s������q�{��$�����I,!@�m��#>ZI]ع˳fCN�x��QS��(^���`X��̇�X衑3�c�~4|�uyx��EʏE�����M�E�z:������3+U�C�� �4ca�ݻ"�E�H%lF�nfr��������H6�}����Pۗ�y�
��y��1��B�fW{��δ��ʩ�J��X/�W�٥6��&�[3�I�`7�;�t�Ye��3��|�18��Z�o~]a�#�>���T�?H>ɂRU���1sN��oB�S.�ߊ5�%'�����ig��G��`)��A�����4*^��4�aw��+t��hAr#V&N�C!��U}�٬N��#������m��0�#a��:�so��,����"�ͦ2ݜ�;����R�t�(�W����G�#���%r.C2��X?�x`��^8��C���f�U,���h7��ÿc�(h��m��S��ŏ�]5Wr��;^+|�{!��#< �jE�E��0��+u����3ȁi��W��>� ��Q�zM���g[Pn���y��Ϫ�K{PJ�k#�$��P?�ZVU�J�k�8��-Ⴡ3�7��Q�/����n�7�P�ˣ����c3?Y��D�Ö,��^s���a8���O:�nP��Z��+E�F'�F����/D���5�'�������)'x���� ���?�텡��HۦMɗАu1խ8;�{mM�v����\�	2]��I��Y)g(a�^�N���k��9�k��!�Sge�%�%0��E+k~%��㱛�ņ&��33�����\�����ߜD9I�vZ���h�d���^؎
���1
i��y�!"k��X-t�'��?�Qr��MU8�B�]���X�J��G~SHo0�j�<���͆���M!��}pn"�І���;��yճHz���:#s�ҽg�2�:��|	��Qw���_����|�E���6����5��|���TP�GP�9` {�s6�計y*	�U&��$�O���9���B�qO���mA�T
J3�ܷ�\,�!��%�ó!M$�d�c�Ӏү�>��bS>(j��$��%S������e���~i�A��$X�����p�T�)�묋�v0R�~e��
۶�I]fΐ��	��Rѹ[3�}K�����{#Ӥ�`�����T������
O`T���ݣ,>�6g�o�����1^}!O�h%�+�
�W�bkdf�I�=�r��(s$�074-�ut�q��q�`n�_�..�bӴ�+-34¨�0���5ON�����K	�y�������� �w(�1y�yDx�~ z���}���@�u~��jWk˕$ ��@Ϸ�v�d*�ԑ�"�!O��"�����=զ�p�SLaZko<��W�hI�GGkr�%L4�F�}Ȁ�.a!�s"PnZSr�oZtade`�����O)բ�X���KS����)�g:
��"���C1�T���Jcv���RT�û+�G�?�"v��x��HZ�ގ�� @����eH>	��	�p��y,Ȫ���Z4�&�/��z9�
��9�U0�x��IB/�f�
�Z\��K$0Y6�f���~1�9�Ij�E�!Of�T ���3d�7���Ś!���J��;hٌi���y��g6G�A��G�=�@�J4lW,�3;�p��T��I��_P�/e�+�IO�D������r�q���Ѐ��3��^��<�ڴ);+y���V`�0�
2O7�g���1��4��k�|���n���� ��{�ǌ*J<b�ݯȈ�Ln��z���q3�#y˾�r�&=���Z�4��F����iiB4���ċ��D#����:�d�R5�`�'��ib�&Ղ翆\����Sѯ���"��ՔP20��:7B���B� �_='Wt�K"��V��
TϋIvp�Q���2Xy@�>�*x�* �?"R�~U'a�.�^�W=�<D�XO9��������}֭�P(x�*8ı"^����mN1��O�|(�$v��4؜3x91jPw��V�*�4���2[��Ql���T��Z�~�@�
�����[T|Lu�_d@�2��5�Dҷo�מ~B�P*�:2r?4MJ�gT���6ī�غ3S��sƯ�8ڴ�,����jE��bXW�[�ѭH�T�ǡo�5��?���,����qǲ���"�8w�$t��8�{ !�Ʊw���ғ8Y�.�8���&<|V�4Û�%��.���9�a=�1�Q=c�_A�÷�,�@x��_!1c��w=�*X��'Έ$��1��x�G,��ؕ0�V���Nه�,bЍ���ڔ]G\a	s���vL�nޔ����=(����O���ꍦ�� �k)��σ4<��$8FHI��IH%��F���;�t��Wۋ<�\�d��x-HF]���M�91(�-�Z b,� G�YVŏ���F~כ��t�z�X�?�0��υU��z�O�BA���s�N"Z�ېΤ��6�{-�Clnt��1!��_���"����fG֕�Cy&���E��H�4;-�1e���Y�
	 +ܺ��Rl�m��P���h�D��ӤO�X�h8%�q�ca�_v��d ��0�N:ߙ��COrd� w�_OS,á�X@�2˾ʔ�/��nż�}"������/!?���PѦ�T�uB�c'ɤ�v����P� q"]b��?=nCD��Ԑ�Q�d�������@��XL{Ԏ�o��8/k4;�`�%���������?x��&8�=�)@���I#?��C�Y��~��*s�,eZ�������n�ƶ:d��.dlZ~[��5����c�.s7���9��ӕY?-l�-����ْ���nT8rjFJS���`iN��㭹���-��V���;�����i���ު��ᑕ;�ѻ���o.��3�3��Mε�r7f��'�pi�թ	�����OiQ��E�)��k��e� � 6Ӆ?��h���1�^C��P�g4�ҫ��!M-�֌����S�k��F�x0S��Rd�U�-��N�fw1^(���P'i­�����%�z�lLƒ�%��c�����=�4��ݠP�5���N�2��=���$����`n���!]�̷*�%pY�|�4Or�@SJ�J-I{�\Q��&�Ϫ�� �0՗;���#6�������>ѡ�n1ۤ,�y���b�n�N�=��������j90'�Z3�m�9����o-9�Z��B+.�gZ�4R(��4�"X���D�*�k��6��y�hP͛2�X.W��T\ɃU�/���'��H;T*� _��Zj(žA��X�K@��[�f�,��%R��,<�P����9�Q� �׻�/߅���s_��x��(�c@�6n�<VC�J��GaH�G�S�l�Q&��d%�xH��*
�R�&WDXs��3AJ��9���P��"��OQ�zER�+MVC�eK�>�v���!�m�h-6o e���&����
H�X/2Z�To��M�i��q!^H#���f#^����@�,��0[��G�:���RP2X$e�I>碑lj��0!T�C�K߲f��1��i4`y-�-Q[sr��v���@س䴏˫u���>�|����<��D��㸁ی���'�я�X��#��W6�o`����u�Id1�l8�9���O(���طu
�׳yA�\��v�z���斤�;��	X�"�eQ� n�$�O�^���)��x@d�c�f��Y�4'	;w�dD+{�������`�L�G7���d����aO0�����<����iL�̪j��A�њ��%�����<�[����R[5�I7� �{��?�л��=��N��Ү������|�̭���c���G�\������S඼�$�/1�/�~��5?� 4�tr��G�W��x�Nsf�$�R_�����m6Ȍ�Ev4�uȚF�jXZ�ُX0=g����Hɛ��J��s��c� �8��O�8��Iul��iJW�o���>X�p�r�lb�K���(;��}&T���ބ�9$W㽔
��d���2"�J]7����!
���f�{4�ƨ�\@璯2���ח����M�k����Җ^5�N�\��Yęq��@lM���`9 �!�0E�Χn�d��u�l/ץ�g�=�!�Q�ג�P3�?�E}���?���+j�R�ƪ򷞓@t���I *��R���)��9Yt���7�E�`w~�Ao;AN�>Ϊ��q��Q��m��E��m0��Б��Х�>��s��t����ϣ�������ֽc���z
�Ke��t���/!?�����ȧ��C�e|�R����}L�S�>6�0p}�������hw���wObK�
��z�sQRf2^�����a�j�T��VH
#����7nt�������c� ��͕>m�3e}@4��޾#7�\��+�Ҙ�1.O��S����� �s��ҕX��D����r�1�� #��?��
�����?<t�2[����N+H�>&�^���qo#��兮j������f �F�v�����s#�:�w���-�����p��""�Z��Mh�s�|H�P`��Is�C���S��sf��S�go���:�06�/L�
���r���Y��^���Cl�\��q�܆_jHܪ|��u;\iL�g���~w�3��=
"�ōf>?~�3���k��x�ŉ���X������"�K�h%��D2[�&�h?*QoI-��;�����0��v�|� ���FH��!݈��C7������p?��'���@���Bz�Oh
-�E��b(�Ie�<������,2ފ�_�
;�gA>)��X|P��-�YZnZDq�������`�@��췆`��0�0�=c���5�϶�>��C}'�ED����M����D��V>kIC�>���3訴xw�U0�u�+�_}�A��W���Q��R��#Z�S��+�Z����EHS�3���3��'}K�u�ߧC�������/t�l��w�������~Ƈ�J(X	�o�^�'g�ufQ�}�����<�MZ�f�ju�`0�ѯ�?�|#!$�~ɓ��§�]���t�ģ�~�4���R�l�Pi�B5��H�q�yV��d#�e� ����L�"^l�(5(~��~Bw����ͅ�䋷œn]�D<��� Ht ^�Rf�P�3i;��2���x�q����pw�$}�L�:�p����+<�h�[X�*l�GE����>�Ѝ�X���C��i�0��u>��7}yLv��i�>�Ѣ} 9S������=-W8Թ�b�0�(�դ� ���/#��b6bT�![�EIv2�터�Pޏ_�����q����P æ|y��oyK�h�ȇ_�D�4����E�	`�Kf�+]��uL����CHZ��:��XO�[��q/�xI�E�3���.��2�o��i�0�r�Ot犢1�~H|�(�ړ0���7���H�ːTd�t�����������X&2H����JдC��!�Vm�H��B�4��c0����wZ�WvU�%RW2�
�6���Z�E�W��[�UVٕ�Ʈa�O�"�Rc��F��_�rZ��Me�-+�d�1��Bt��O���������v�3,�۹I��VҖ�`��|J�����ė�#|�p�i/���p01���U+���i��ԋ��;)��=���-GF������ޯɗ[e��*��0����TE�r.b��{�d��7Q$I!]R%�J������F`=x����N3�{�,��84�C�S��q2�ɠ�y�,�91�<4��~V5����_�z侲�d%�1��.�}�Q���lh�Z��,�:Vd�,�l���gI�W�s�y��������TH�g��J�-�T7�� �����v�x��/lJw1h��cAhI!����úe�u�?�d`��?��Fo���wX����9so>-N�BS�xK����1᜙���5uٯ`N�p26��@dXg}�*��|��-E��YA�	�z�Ü�!2�)��r�DD\�)�S|�J�$&��FQ�	-d?��xEuM�̀&��bh�����ǈb�� ��F{��q-�Eu},�=���S����#��N(�'����ޱz:�ۅ9؈�?�n]?="j�_A��?>F��b3
����Q9qmvT(ц��d-l5�������b��k�� �<�b��0��������$g�8_��XV��p���]��.�R��1K�1�(����c�M.0��I�����f��f ̬8����O����n��3\�b����hB������
ܿ-Lɪ��0���	̩يS�w�h-���yA�7Nh�����=���c�J��@X�0��UNB�C1"���12FС6����U���J��|{7o������E0t������NU�� ����%���y<���N�-�ZT�hǝT�x�<�6sb\��H=_*����(n���"C������q3� �����t'#ŷ�f-�N�D�Φ]5�x]no�������i��s��G�*O�S`�w��U��
�r����E�\�嘗>���Ň�u]��W�P�so|�IC�P�Q�n-�I&k�J�c��C��F]W�i�^1�v�� :� �ZD8��C_X���A��6g=�b�ñ�t�	/�4.F��|�Ͼ�Yt*��du�ۋ��|�A�}��K���Vcp�@���`�Z�%����dV!\�fG=�1TG�yr� �.wkY�"�a6PJ��&��g�!,�)�!�� a�eD�f��ĳ�el������ل�M�]j4��f�r��x�0����K���U��aY����Ryh�ܘ��%0��t��ćU�D��|�QDHd�s������<��Gp���3�9���-I��Y��ώ��;�~F��R���^�ZC4|�C�Vs���1g�]w���8�\+w����t���~L������*��+Q�oZ�-�����Ph������0!Z�-CJ&
Y�ty~��6���LQQ?�C��En[- :Nqq+�#�/ˎ�2���̷X��eױ�ŤsPVu�)P���e�-iy�y��A�B�^NK%��>P�X�+\g�u^!`�i^~����)V�U�טmW�	�qn��p��Xr�j6�]q^BO�5������
����Y�� L/�%��;ĸ�u7p�Vdr�E"���w#�gq�[E�o��8�@���<�g��z�u�*�L�T�-�خ���Ƥv=W�a4:'(�EN�f�*²���M!�K�Oa�M�I��^�+;����ӱ���Dg:�i��yKA���23�+A� }������@:-
{���_�Nvnz��-�[r�e���7Drj&5��ں�zȅl��8��'��R�q�Yp��)�nD>��f�PY����,~J��[�0�d�')������Ǎ�U�1>&R|�ow�QW������ "�i�>b�C�9)q̩�Es�����%�9�"�i�34	 ����_!:���ш�vp9�s��ş�孼�� Q��-��?r8�cvݻc$���I䷐�&���|),��tC�� _Z��G�	f4�f�e��aE�]kէ]'$�Ӳ�1H���`Zn�Ԟ*~��'e�Fn��:��Z]�S0v��	]=[�6��3x."�{�� ��Q΂���Ͼ�3	��w�_�ASf��!�eK.3��|�g�M�X��WN9k.�В�NZf�A��׋�,��	0l}��7r���֩y��"�{��')R�n���"Q������a�S�5}�����Wk-��S���?%�݊3l��ۯ� ���7�,,j�����T�j�oᝈ��	ֆ��hŘ0@Ti���=�F�_�L�iU��#�(L�v׿ZNB[s�VH�l�>!C���b�;Edg����0oZ^tQ���HK�J�C68���C��������>�쏥:��y��S���l�+^ /�]=�Rq��y� *Ez}��W2F����iAQN;5�@W.��c�� �fߤ�^����l�+j�k����-uE��ߊp��Z��0_x+-�T\5�O���*�6��!꾰`C5<��*T�	k��Q.�;P�M�K/�8��j�X�=���I���Ϫ�!Ib��]t1��	H?6FfW������0v�oM|ʕ���%q>T��c5�#��C.1UX��ݴ��o%�*��/1*4�F��� ���?Y&�B4����]���UM��N1����I`�?��bqq>�{�d=�o�P혳>��Ogc������t�\�dl�_�:��zo���T�K��I`��E�F���מ�������S�� ,W��u)]��8�V��J�� ��O&���.=`�\�s��C��Ƚ_��jd�"��s-<|J,�yEݹ궠���}�ֲ������l_�9R-%Q����l�������UC�v���+em��Cs��S��,&=+���:1��#ɭ�Р|��o�E�!�t���pL���hs�a����dq�s_�5m��7tKsҒ�z�5���>�l�`�YDf_#XB�f�ysl��g��e�ܨj|@DJF��mN� Ԕ)4�5�(�˾�>Xtޜ�G�	o婌���2'e��ϑ�=����<�y��4E�ɺ釦�˲��gd�E��l���h_��*��Ss���K)q!��ޡ7曇j3�{*O`�@� ����؄����Y�N�1s�2x��?�܂|[������k9���*0���e]C��7�L��bMT���nn�R�Be�����7<�V� ��j��1�9�;2��}<}�C&[e��7�u92+�pM¨�c�e�Q�H��'��H ��_z�7�٫vy�}_�%��9l���{��ֽ���1�T��O�c�s�7&��=Yw]�%l��;�?�������.���f�\)vȥĄ~95�t����Z{P�$�:5�V�i<!�� ?�pH���R�ؽ�RW��_�M�}h��s��KK�0��G�砾����>b+���]J��ƚ�P@m�=�`|�m�o������,I��c������lt�$P��H���;�p	�߆#s�*�B�~��������tF��f¨L�A�z9Uݦ�L���޵ �rE|���4�8'ͧw~-<T:�*\��.@�,g��F� ;D�5)�7���g�*��D�6D�C�����)rΞ�Z9�9�Ж��T�tH{v�����8B��uGںq���S�<�-F;��m!M6i����o�?�Z�1�c`a�i���}���~*�$)�[��3�$? W|�b;��>�(�Y�ϺR�cv-D�Ʃ�u��L2B�4�&�5n&�.���n��Ⱦ�J�&k���t��������S Cp�o��h�;*�Ƙ��Z��R��QI�	z,$,(��@{��JCQ��@>:l��u,v����u3?>�0	[>Y��5DW%kU�߀�wG|��4���lr���6�,4��]��A�db�%����s=��7�L]�z!�Fj�-ť�F~T�]S�8��3S,uB�zW��\P��~�RYkM�0��,}�oy�/=���(��X�!J��t�3�7n��a�;�t��b�Z�����h��+��W�-Oal�j՗j��X�.���^ϭ51O4e��,��jN�"@ �z���7��Wv>��s�W����#~}���JR��8�`0m�HQ<óIG�/�aGJ(�d2���!�\1���u�ǆ��j�Ȋm���f��!YÿD�����!x�'�}���̼� ����[��8�����h�����8�8�J�$��r3�n�8��k#��@t)''wp��p��l�UxQ��c��U9zw��JU�����l�К킗3d·I=�$��b�s�������]��5ĘjP./?��[5�^+w�@���!�g'I�sA� �b�5�����㒕[�m@��|�m�:8�*#�v�ˮ�U+Ê����sT�jLD$������ѩw��	���:x�2�*T�;v���q�1@�(�j�1�*�O3�#���u]AL�*�̗�Y�ZM>Ks����'�Z	�{*��Vۮ���OB �Z���7J9���ѱ|�]�l	�G���R�`]\	�l͊�0q]������%2]n7��3�:!1�+z9#I/�1~U�IU��u���L�0[���y���ȓ�=m��� �)��=�D"7����F�J=��$M�*�0N �Xo6(ɻ�眸�����¯�ھȦ��m�Q�z,��ڷ���|"�J �\o�D�;ui��>�*f;� ��\)	v���_R�<?��Qv철����-��#���8{	�+q�KY���]��d?1d����s\��<��lA-���������f�^Jd��q'���#)���6��j���D���a��G}4���6�7���XH'�+�lqy�p��f��}�qN���ճG��d��E �L��T+Б?}�L�X�n���U���E��ݫ���Z6%��ʉ7Ee;#W�R���� �����:�x��2��,d?o=�M��Wi`�P�q��/��_��J��eQ���Z076ʨ2�r�~Lr�Q%.��_��єP\�QD�i���D��1U���t���68_s��|{sod6zr\�C���+���14̓�4O��d��z�t4Ξ��d�K�I�d'�F�����G� ��>�`��e��V��|�k�5tY�1%M�f�Jp�`9�q�f��M�.�ؐ��ѭ�m:�?�G��%����.]����f�4��!�=QgSj^�Z���dY &��2�K��}d]X�**��/���� H��hE�M�Y�=��4UM).݀e��Y�%v������Z�}Y���5�iϐ�|]�ʝ��lp�	��o$o�� K�Ι��AՒ���Q��A@|��\�c��$��9R�I��u}?�vi �P��bkq�����_3���F,��B9E�3�7�6��lc}��x2Q��V"����M���?�A/t�_ԭ�φ��qϜ�,29t�8y\�O؉�rc�  p�C8�jxDsެle|/���>�L�pU���D��_w�}V��&ݕ��@"���,�%�Ԓ������~�x��5	-���ة&���?\�D���e�BO����D+�c�M�>�R�-������?$l;�+�ϋY�#Hx�W]c�O+���V�ӵ���X��(&K����n!P1l�b|O-��c�"~p=#�#;/m�`x�BL�M����ʜ�� �M���_�]�&#�Gè9���KP�d^���x )��&� PN!��������JV;���ʳ�(�<���S�5[GG;�B̽��7E��N�D�.J9v�(���L�Au��>_x?&�,�&��O�G��2�H�r���T�-�	
)7�2h<��ձo{R������;f�QQ�B&���X�,L}M�����������B? FW��F{�U���J%�Z��B��AB�GƖ���k�Eez�:߮�5Dk�2"��%�[D�,��e�*]�$ל/��Jq(�p|��]�Q~�_�)L�z�8M�k�kDM��[��������^�m-INa�a���Ӱ^#�D^;-aĊ0�� �W�cT�'m:�*Z�T)�C�M���/QT��������]��y���bݮ%8��6RE�e��a���64!J`{=���
ۀַ(Z#������n[׶��X��j�M�'�xTed"s`+����!2/��y���张�
�k�[/�K�O��l��N%��,�a�̊5����y�R�	��L���c��\�P�!�#"j��$;S�1.Xl{<���%�U?�;omw��!������<��&�}�x5�
�~�1wW9#�>7�w���RG�m�hv65�ЇK1�/7n^9�U�aY*����E�DҒ��Q,	fv& �ϔJ��y��J�@���ut#��h:v~Dͥ��9��R�}N?E��v��6�w��45����vָ�7�pJ����*�c$�VwQm��Q# ������/��#���,�
�4K�K���^�[�D�*6���P��nԼ����zdg��҅�I+1l)/#�cJUlm1 qC��廋�f����9V�k��}(���C���s[e1K�g�^(�>Q�?�0�*T��)�a$���:k{s�l�ȕ$�]��K����W��5,*N� �䀃��1�,��XȦ�=��kR� W,�t���Sи�%�/Ӝ�s��X�(�:�UƉj��o&�ſ�ݱ��#��ޣ��W"�ꍁl����j_Sz��r�2�=~��<�U��-2��Ԯ_��i��-��,��b�L��4� ���~I�U����V�|s �+fK�������E�98F|���#ĮJ�_��d܇Zw�(E$ŭi*���Fe����1��u#�8�I�GB�3R��z&�Gl�{8�N���h�s����_��j�~W�r?<�{�+goYH����zU�.��	�	:h��R[W�d�7�XP��K�TT�d����}Q3��Z����Ф�����_M�eY�n~�>���7y�`�`�DD�٪�^O��d�9�kD��g��\x�r�493)ڔ�}Sr�0��y�,��`���t۔	Lk¹X���M���t�q�^���dy	�Z`�GZ��o���rB���"|{j�wl�/),�wH"��r#Cl�W�r�����<6�����w���y���W#�f��΃#�ˣ��iGD��u��$���Ix	�4��P��A���F��D�p���{$�a3aj�o+���T\��l.�7!0Wp4o���}f���ekn�����]�,���`���ڔ���J�` �LK�ww;�.�0:M�I;b~;F|�Uƅ|l�)�y�x��t�k��+��_�	@��8���ޘ*����T!����X,���.�WT�I
�MS:0I�҅��D�j5�-�*X ���U�����;\tA�8`�������8�BB�5}�i4Gz)[�M����^7@�{�?��P�ϥ����,7�ȟdFMビ�8�}K'�B����T2߅�d*���BG\��dL9�$�7?
j!Xk��=�$�p.ع4H�	M#�
�&n��s7X.��OXr��Q�P~l��z�\��B��J>٨�
{�k�=J9�5���"�����m�I��(ߵ���Q�VHSq�&W��V ����d�L�6T�tD�*;��ƽ��}�L'V���[X�Hʪ��~u�5:\����מ��_m'j�HD��Xsr�Pg��9�������5�����/q1��ڻ����
��̷�b�.�	x�13G܉D�Ll�[U��3���M@Wy���%E@ݒyu[�^�t�Ď2��M�y�%$�*��Ϙ�I��>����@��}�+U\��.��F�a��B�O�b�[��G�ڂ���2mn�+U*���=G��9��9Ϸ�N��qY�;�!>�-6�h5+�M �of~���gY�J�@Ȏ+ދ�樯|	k����<J��nr�(u�o{YlR�ew5t���$x"�X��ްg�a�?����8��s���7G�/Z��j0����J�D���/GW|)/@��O���8,�*������QS}f�*��j4X謾�ߪ��|]�޲ T�QxX�[�������F	ĭN��T����,��������y<9-�`,H�p����E�,�nT�E�ĥr^�(������t��8��:����XB-��W�B�NM�!gB�C��}�}��%�Q�\"���_��2�8��.�R��iw��_!�8��+�T�Q�/�;�����?��b��D����Յ� CK�Kk��A�!"�N��Wi�J�NI��#�%�I��2`�	&O��m��H*%�f�t�*�Q�p��Z9D^\T���V�VL��Ų(?�fh�yؐD���[�e�nyL�K�ԟя���r����(�0��?�F��T�l\��Z6] Z.��"��?��M8&�W��
f�h�1Ĭ�����*���~ZH�@��o�.�����`� �y��m�ȇ��;�ٷY0�IU{��
�<��#`Ұ�p�|<[`�+�_�b�~��7��l��beW;��u�?�[x�;�2z�>Jr�h3�^?���RB��|�-m����M�D~6���2	};/\ؖ�əS��ȅa;���;(�\6"^�ډ�H]��a@O��
R��F|�N���g��f�uv*�B��g�� ����Cͱ'��u|�y�oF�x��YzW�n��A�E�d�\��'��U�<��N�"I���3)q�P3�@6�7d`��q�qY"Wxi�� � �r}DFym�Ĕ?<�J��Ni�x�ix������7��_��i���Bu���镇T�����F+���#��Tİ��hS6�� ��r��?�%�Y����I�%��/��S�<��&�"ˑ�5�I$����������i��*'��m�̰�*�����i�jO�ypS*����K/�����ૅ���q�xd��o���!\��#�q0��ELB�nNt�QA�� �+&�FP��	��GtT����SD��\f{=��p��ƪf������Jv��q��
�]�������Z���eS#)o���b,�P@w��g��k���"������$�sCƟ�?�K{���x���i/i�������Ѵ=+��uc�&�(��}�b��'ֵ�4Ϣ{2;+�e?&I������NI��f ��5@�O��N+B�MiP��(tP�%�\�Ni��	j��aT�������Ѿ������u�0k�R#��pmF�A��'`d��_�K��19��1�!�A�<5�!\�7�v�!�LBq�����Ҥ�9�D�[���'O�?F��D����&ݤM-7"��d���Q�}�w@��f�-l�;�
�h�}��G /o�`	o3]�>��������j�P�m��್i|����p��9켂I<b��CQ��b�p��Z3��05ˆZ!�4���'��6HG��]x��������xb*i+j�� p~��tۥ>V�i1U�:ZP�g �b-����(C��\��֓^V+��YE�-�Ԩ���"�8�g��v��v�n��;��A
1"��b'+f ��/;̨Q�u�L����E�r��i���d51������n~6��c}?d,m b�K��*��r�Br�RZ��t��+|kPWkLb��%�tn&�G�����F:uv,O&?�o�����7�1_���=�o1f�# ��ѠZ	��s\��o4�>�Sl�����2�$?���"&mt�+���������Nyɽ����وJ�1�1���ğ�_��+E��^i�!
{�!t�!d'1,&������&P�<�Zyw�Gk7�Wќe��a�kw���iw����� �_�����
йtr�0�)v��6��P�)q<*\�,��s�\�%S�#��}H��z��ȹ�,E��w�]��@J̰�U{]��U��?[$������ۦ����V3�,Q��=.�ֈx�D�'m����^�8�!��'�I�87*�>�g{DȂ��qžk�v�7��Y-}ie���5P^���I��V����ڝ��j<�3u�3O��Q4�}y�w}{>o4K�\�_�ɞL�sU%�{iC�ťac�P�ա]T��Mܗt������u	���g�3N�T0W��1�3)=Wl�q+�	���3�.5�e$������= �\h)�>Ix��љ0>��2J��wh���;�-� ����f�j��lTՓP���� �����T��8􀈦
�"�J�,;��O���{����(Dp}��]ڬy����y��N�P�摜�n�p����S2V��Ɗ��2Z̰�רx���z�"È���s��8=�����!q�n��u*�"I[�f_kv��L�;�^w��g�l|c����IV:d��[lX\�O �m%��Z_6��4,b֏�E��#U�G��,#�"�]����ՓjVh��z��I��ܿ�U�+�`VJi�N�4c.	ϗ���wmX)E���D{���\�(�0�OԠv�h�h|��
nu=ݕ�vp����ְf7�L�w��Ͷ�.ܽ�n������o(�hg3bq�1��z��iS���Wj00���hF���=�YV7�ꉍ&��h�k�32��8qkd���X�v�M#
���LL���q�[��RSp�n�D���>�q�A���K�2��ǔ����L�j5JOآ�
�&s���[$l��ٟ���
��Z��)���Ҙv���v���D�.�0������������q��Q3���ĘL̟�$Epo+ J'���T%6��A�,�S��̧V{ ������ⅡUJ�B_A��kW@M�S�`���n#�&�uiW�c�J�}�x��8<[~W��P!G^���E �"l1��7q����a�.�L -��I�^徨5(XK��w� ��U��'n�����ٳ�+8�e�!�)`T��� �G5u��F��
�T�m�	7�π�p����{�ڬ;��݉a�4_�x֩�%��\w��>�Қбb���]c����|��A�~�y	D�L>��Gp�d��H��K`��6������.�yXW�5Տ���f��l%3.|�.a%����xC��W�m�lX�˓N$�6��RigT�M�{az���k�q�$��k�5~p��R�2�D�.��8�c
�,"5���^�|;�={[_{-Oz�įNϑ�{v?ά�#G�Q[���N��[ ��'b��J�;�3�����9�����F�Cve .��o��w�w�AK����^97��8����q��\��P�~��U��YB#n��{pN4J��Do*k�:>z�}Gɥ
��e*Gx���V�
�����3-ur�S鳽�5����P��֝RKQ�e�ࠄ*
ڣ_qA� ���o�bEʚ��R#w g>j��ny�Fs���Y��}�$򹛩�ҠG��{�P����Ss^AI'O�b�4��$	����Ţ����:xY�h���>�GUvћ�W~���Ŵ���K�I
�5,Y��T�7NJE����2="5�佻���$:�=���퀘���w�Yr�)5y¼B7�G���� �P~�ݥ���S���5X�:qB����J�
�����H�WRR��w<�(���)ҕᇉ�?v�}>4u�E��[@G�Y��f�(V��S�i��v��ht�E�}0q@�j���4!Q}�����</eL�g����=�|!Bc�@�כC���!#=��в,6z���|,;�y\h �+FI���T�����'��z��s8�7�Q�K�F�2�5��a�N0��vI%�z�?am4nP��o`����g��I|tVS��f���j�X5�O���ђRӣu<E���k6
��U����^��?�pCp�ӴE���2��ﳂf�)ݟ��k�/�����֨v�UBf�ר���b�� G��`�[G���)v�@$8iz��u�4�YtD�'��&�UDE��Zm��NB�+й1����w�חn"��a��p�6Fv��S(I�J�`�A��:g�ps3\�˟Q�0�.���z���G_�j��:I�ٷ��2
�J`��B!��Uw�����8E��A](K���,�;eٺS{���L�`�{��_pg���-������S�Y�-����<��ګ��>�Zфk��H�;���Il�����(��k}j�w�������FU63��BQ1)f1��sOS'��E�+��A���(�%�x�/�F,��՘�P�鷽w�/>Yz�a	ٌ��{��dmޮs����M[�m+���q֐.��|c�%���dS�1�l����i���J�D����n���w�=|�	}$�yg%��t�p9�	��ڪ����
[k�R"f�:]8�KC�`LW9�g�v}�X'#�j��U��Fq_o�5��YNj�gO�Ƥ�R�A��
T��,l��?�!��v��U�=�#���BT��h�Ъ9�̕5Y>v>[.j|`��%�̜	���I�Z��HO�+��GKi���'�����7jN�c�]��\H���<�tR���SXr�rO��>����ֱG��A��k�&���h�>��\Z6��}�%r���~�L�r�_5�^��n�#L=�0\��+��g����iA((t�����@�E	�Bձ��ʦ��b�Z<���N�cEQW ^Q���0�ۚؽi�9>��@��3_��7� 2-򘶺q'dhީ'�Ks�$�)c��k���/'�l�1��d��Fڨ�j(5�~��^,{�
#�.3����f�3~�|k�oR	=A4��%���~e$�gs� G[�mT�B��x�g�a�­67hu�[v��#N�Ki�@�Pˌ����UspL;]�e3} w��r�<*�=Ae.�7�D�G)�*��b羫�WU��ݢͿVYr��*i4���Ѩd}�?~��������?6���t��j�a���@�����itw$�|�W~ݰd�J1���E�	N�����,g���B�tÖ�/+��׉(P��� L@�n�M�W�i���>=ԡ�(����+�k �8�Q]:)��nP���S4�*�1Uj?�h2���e!�
i��$z:���p>X
�����Z��(V/W*��E~5��dk����刅5�=�v'�t���u�N��"֛TI
��;�C#��}�L��uy��*��Fa���p��U�?#D���O�S���l��R��08��B�[��T�[U.?9{��F�ȂEۯ���Y\��g��m�IΥ���ѳN�넫��P�M������`�8HJ�V��[��6�>�A-ȏ����@{��%�S��3�'Ҷ�a_�����Jt����6�vͪ�+�k����E�GP�r���O�ws_��q���%Sw0Ք��_|�gѳ �o%�i�Dъ���+�{E�&�ÅtZܡo��9G���i�� �<<�Lt��]x��:�.z��>�j�7��HwN��\K-Ȕ�|@6F�Ϙ���֕�ԁR�t(��`�:6pR�jo.�}���-T�>��xq�6�_�߆�֨:�S)"�f%�v�T^z��B��?����q��	jAa�vC�	�Z�AUQs����!���
HK�����n�
�+��� HUD�Ԋ{:���~���R("(��mIr��L!�0U�u9 ��M
��k\�t�W�$��8��:>�ވd�n}�_�y~N�zT�ȗ{����g����F�U���}�e�� p.��0�KkR̐��^I�B-���M��F��A�S�vB,��:Q�b�	7�#~�gLm�+��Ձy,Ơ��4�p1a̾`W��K�블Ue�yɨ(K����>H��#4�ӡ!���.�)A� O���qu̬�W��~��PN�Hc�z���2����wq$�dy{z��a�z�]y�G}��RL	1O�����(. ��U[�צ��n"G	�SU�5EzP�'�6ULJ����m�䛦�[B��܇ -5t��`[QpƲ��\�G��c�i�|�&>�����R=���ƷJ��y�+����4�0�Yv��R�l�#t b��ܪ�V�hb�?�]L�UtN�h|�I���;6a6�xx8�A9�]����N�v�Qu�;%�Hn0q������[����Ѳ���ʖ�-ǂ{�j�f�(�e�LSwOO�}��z�#���(G>5��l�Σ2k�(�Ź}?qP���6#o?r�n��3�D���9��C��+�{�w���.2�J�zm��O�Q�J�a�%��Fu��-(	?g(��t�|M3�B�.���`���w �yO옐U��=G~�h��RߦoQ]F����FǦ��C���fft�`��ʣn�Jǳ�۠x�E9+(i���䄋�hw�&Y7q\ٴ��D7�\q���].���DH��#S�H4����IN��:X`TQ��K�7w+v��Ǻ:y�e&� (�ᷦ!4,�F�ռ��W�-Ь��o!�����/ߗ��Bzh���8Sn|�-�F�h�{�+�-�G�h� �@�*aEr�^�ӧ�a�ZD��;^,l�X��>%�E�a�렖��,g������c��\�P5���N-��X�c]E��J�3 $���/�d��ͱFN=-�c�/	{�����x)�[+��O��c�
�
Lp��1�~��U��$f�$��6�]\�q�7��'��l���A[��7U7؁[��X��!��������YQ����l��P�M��_�m4Z�͏P٘��;��8v����,5��;x� p��#����l��?�N�Բ�	� g�h�!��8Du�x�Ŭ��]�G���J���.������"vE��ެ�eoh�P�U����g���b/ �l�WZ=Ϝ��^�tN8�
�á�����0Z@=��>�a[?�4��`�b�D]���{�'%�؀�T;f
�EdnCߊ�>-9��s&){d6��������:x b�|���u�F��Q������G�d����+xb\/t*�t�ZOsx�֝t�k3B���ؠ�>��!:��wt��ɶc���7�kaxjnz%޾L
��� f�}��F�")��I��󿆡e\������ F��l�Wԓ2�"�a��х|T!����wDLu������ց�]Y������*9w������p�H�<:'�{��8Ւo���S#�����y���mʾ�{PI{=k݅輎-*�A��k�j��-P�)M�.��A�&�����@�b2��\͞�2^
�Uk��o�4�[,�Rao��Sw@5�;����;��dA��������2;D�J��'X�VY�����q�dl$��|}J�S��͌�B�׀3:d�/%U�(J6��y3��u��1-�x�"����'RfCqa+�<�[���.���R��m�cq^Z���+�y�=|�	z���Fg�I-3����z��_��h�����S�vb~�!?�Dh1i��!�k d�7�����M��=N��v��d��$�u�z7�Os��KYW�����wG���lz kJU���@[��#�� �FB�*�Y��m_YB=��Ve�=
1�gx������N��U��r�+�cQ����}վB�~u;>��ń<G�f���3���+����������P��D�����>��(y�����Å��Z�5��q�����z_��&��4>~�l�hW���~�{�����N���|�N�₟��>0�]�9�t��pZ�O${�S��yY�� ��N��MC{�)vʫ�8�!��nYz�q��݈�ǽO�lw�� �g�i1�_*�����z��p̃�����L�FUi~*�0T2�:((��!�y��º;�G�=���(,e���8��4�0�3��&�\��z�X]땽�K���S:d���M7~��p��%+�7Ζ���5�iƴ�*����B�bbn4Jn�Z�g�`� �cy�I�'���]�K��:��4?�U��M.ձ�*��~|G]W�ed��<�[3{�T��	&8���L��)P��?���k�X�V79�[�̔b/F��Яޒ�� <��'��т3sO@!A����o�G.ɮ�O)t��УW'd�FmF-m���o�o
����6��-�AU�L��È�����f��]��9��G5���r|z��I}&L"���HiL�P� }�37m\��x��M��ꕖř�)�3���pLnG�9��Fc-Z�n4膫��c&?��i�_���N�s��.��ü�cSm�����I�o���%H��P��( +���I�������+V���SeE<�~�1�q�3��>�T�6�ٺ��3ʚ����Uj�!����y��1J<C���/!����OE�V�_1�Θ���Z���712hV:F��-���a�����GȫOݐm�yٶ�_�Jx9��;h��k߰�|#O�W9!W|X]V* ����[�QL�Az���3��F��qX.�$��`�G�j\<ka����
?]�֩͸TM��Z4c*�Zz���c:��w������5d��c����V��f�N�|��%��k��l�m~��*4 K'Ź@�M�>.h�hҪ'�ш�W�Ɇc�
�8�L,>����V��x�զ*o_�[��;��Y/���u!v�O�od���cEǚ�
P����������S�����"�}2�C(��>�z��G	��"���i<��Q�����Kyp7X�0�qN�f��%i�zg�=���C��V����0����3�@�%O���h)lI�ϕQ+eU��O�� �����/\5��Y��O,��sj+��Wm�&F��~���]I-�_V��$ ��:k<lJ�����,���R��E����>V~	�y����i~p�s���:�Sҏ9d�I1ѐ:��r�Z�`�/^W�q��ģ��'%f�cF�=𥊤�� $N;j���^��%b�Q�@=�0B�+��ޔ�1�&�.���
�����#�$�j�5)
7sBf:�J�!�X�'�Z!*�ܡ�bZq����k]��`��立�
�&���oTy�t)-�5�A���9���8�V�����PؐiY�!-
��(F�UOyC<�lpE��Ȭ9�f)Hnb�=~cr-��6����~בf�X���Τp���u.i��t	�e�~j'�G�}
/��K%��mLN�F����kNhl��͙�Z�#HZjI{�G�\�j�� �K����O҂�2y, 4^���f�ի��{����l]�y��d�W�\ģ���n��qY��D8ThǥIS�2c����B=.�T���M��m���D�6�!�T 2�O
���׈r��h��מ�A�G��T�/ #$d::|�Xˢ!������^����,�H���xtU-34�S���4��bG��E|�ke�o���"��d�pn���l{��z��v������5��w�~��5f���8�>�4�E�2��t,�T����ؕ
%� U7��>"�>��Z �ʉn�C/[�Є�[�y�e'+:��Z��_*l.���c$w�:EX�'����$��PX	�>IU�����6�f �q��ש0�9^�Z�i~��E�D�^E��+�riI��ʸ�eê\M��U�E H��w�~�րL*I"=I�M�U��]1w�
�/FqT�C�e�/f[W_,�!��!��OX �M�BR5��V �4��M_/�,PH���~�.��R���{Ü�:7���tis����h��&��(o��s�	�_k��+V��w����=H7_�P�Y�/�K���%:�󗶅�Mkv���z�b4��z�[�K��!�>sz��!��q}�N_�' Z�2��| 'J~T� }q��i�7(�x�7�	�<!kл�"�H�1�}�6t�5�RHSo�&�a�a"/�1�.�}�%EI&]u3BZ�>X�Ծ���O&��q:C-$��,�4(��	��덮^VF��+A(�7��4W�����*�B�g��`��!)5MX�����Ķ�R!�-j����B�7G�u��\�w����1�/ut��v;�e'#t$-���}��Cy:B����);tXD�(m}�8<-%d��F���d���5�Wʧ��~��Z�@(QP�Z,<�3O<c������6]~T��"��X���T�ciq��q��]r��ipRx"=�V@�f���^q�&]�dAzJ�e%�w�S����JƶoA����fr.v�C��̏(Zရd�0�{�y#���F�iF�c��	
	��!
{��b�蹊\�]��BU����)��5�$%���U���^��4(������0���]���9��c�a���#h�z�/3<2�j��>8�"�ω#�n>���'^�?H��fn@�=�B��[m���8��@�\nB@�صz?�W�d%�l�Z�k�?)�qj���%)k�����LEY���T!z'P������*�����9�)�:��J��(M���^�th�<R�p3�j��
<�ׂ����/�kpk���Rs�x3nc�wIqt�;BL=���1v.�,�gm�aP�geAtV�i23xW<22�nm�-+�n�ѹHz8�Ɯ�z�$c��VU;:��)8�ğPm:���jQ��1�]���.��ʂ��n�C*
BD���Z��ʞ�eB�7��R�6��Jİ2��)�l�=ǠW���P��W��]��Tk珷�p�Á�1	B��tu�PF�ܮ)� ��$�&����0��nC��z�
��?���ĭ/%���Fjuʑ܇���}��)	o�s�=����gB����Ik��2[֭�&���Lu�J��4��8�!K����T�4l��ǌ	e�'�@����\o�â���D���=�egxk���
117T�
��ΨO��n����7NB��`ft�o��Tg��@�h ���B\M�7����:RR��'���G�sSu�w�h&)\��U�&��X˗xX�l'Q����_��zX�0<M��zd'�p��E��j!�������Q��GA�	��cu��5&[�����A��g�)�,���q_�7�����6m80F���u/�6R���|�p�(*���gA� ��gPƟ.S��ӖsL��n��'��P�1��M㪾�L�}۔2�$ͨ;��/�Ƈ������c�CFħGN�m��*	��}�)C��M��Kz 󭝳I��N\Ź��	�9{=��`�o���4c�GO�X�J�;9H���&��	-�U� T��-���B�%�sq'Q^�U���V���]��:@��񈤹�RX��7lU����UF�>:L��nOc/rj�9��Q���J�iRZz�&�@z���G$ng���@���-����el�8��b�Θ������[jFg�4���n�}@�mD����._XbM
�W������i��q��/��,+��嵑���R�-qTf\���;�I�tɇ˚3��g�m�A���9��C�z\�~v0ɑ�' T�%�@=�+���l%Ƽ�B�B�R��{���tN�B�DŲ;��N��>7f��,g�EՎ��ʋ#LsMɊ(����f�`1�����B�!8��8t4�PD�VΎ5r���ˑ�����X#��ő�i�Xubo�J�yl`�XYKr�C�G~��
Z>Q��<[@3߻��4�NB&��3��k��E�Ϲ��݇�V?�ö~#4�dm�xzL�b�S9��8a���S4J�u�KnM�M���ɂ�|!^���7�g~���� W&�Cȫ�e{�>��Y���SԾ�GT����M�Z�5Af��S�$��H��_~��!�Wx�dw�q�p��5�騤����:Y���Xz �����a�W�a��4�jU<FQ30����;JL���VL�m�)O��kAG3!U��<Q�Mrsz�}z[	l7���	3rHaY�,���|����w����F#��AS���{̡֝�7e�K���_�= ��A�פ֊�{���	��^����
�8x_�� ?�g���ד��Q�ZD�ه麭�PV����}�� ��_H:P
)Cdg�ю>��m��>�����q6��>O_2#����W~�:�=2��$��Wi�r�I���~t'^6�kmlek��		�ޠk��&�n������g@?.ejI�ݤ���N*4T�I�E �
a����d�0��
A����G�,vى=�#���f4���sq���Ղ�&?^����f�2Bseo�?��ڀ��@�M�����_�L���OK�)��k�Z5�z'߸ֱF��� d߿��[���ѥp�Ѭ(��I�T��"����(����̙8�HQ�0)E����D����YvH�!�Xg�Sb#�q�
��I��9�$�S��E�N���X$�/���+	�C�{�iH_e&�m�e4�*C~��:O�/���PJ�rd]��wg������2d���g6�?�t�^�I���k�i:�ʧ]h�2ɠӡ�!#����=�M8�F9�(�B�����0nɐ3�̈S�ص�Re�����GRܵ�z�}Ǥ�&L�~�A��i�E�K�[4-\��}�O�$:�Y�>�8}����k_e��`���f�}�!x�G��it�gV��sQ�"U���l�������s�Y��������4v�^��^1�T�yi�D���ǰ|�*{�e��zd�{��.O�15a����M�a�4t^ȓ��N��]��vd�s I�肻K�Q���	(�:�<�m�	�Fq_�j�6�!rGck�m �þ�%5�;�e���A��_�PQ��6���L �ɟ`���^�54���d�z~w�K����bk�Pk��@cH�v�v��M��&i>$�)�Px�ێ=U�8STCo'�>���+��L�ޯ&Ƒ~3g�f��H����]�ơ�U󟡢WB�
Ba ���co���y�_�*�C�)�=��J��ChvK������T��\s���T���˟ 5�<2���)�X�ͤ����L���c(m?L��{��,�>���J1�zƇ"��s�-?���>j6e�e�k D:�������C/T8Nv�1�+yc���ͭ.SDǺ����5H,��⒨�$��� �n&�uTwW7��n*4�� �=AI���(��]�Qq��5�������]��hB�v������5��J�}���$D3���Ɲ�i�lmy�3�ތ&ZlV7S�4)ySWҀ�������9�#���4^��X����W�e��c����؇P��P��ǣ we}�Hn���Ū��6�೨��(~\��*�G�;a�NK#���0�忳�W�� ��C���U��0��n�l݄���C��h�6"N뷤=�TFZM���s[��Q�<�"��E�E���#u�����x �k�/
��g�#�W�c�WdF��͋ojS��ľ�!rfǩ�q�I���h:�h]�����EG�x�˷Ӟ�W� ���C��g][i�j|�:,�ܤ!�;٩ΖW����	�L��e\ �p��娸FW���w��B	R����C8�jI�d ��f�	(���K�|K�5��~/!��6��s]sū�P�+r��:�#i��M��Ȅ�x�[����=��ʑ42��;r���!Ҕ�Hs��ܺ�g[k�kn�!�LP��f�K
j��C�vL�c ���u�M�6��?�6�O�[	���<J!���Iֈ��ꚵTA ���On:d'��?>�I冔�P�1���#�x0ý���-E"A򯧜U�Y�i��٤��W�����;�>��D+��8�4
��*�%O~ڼxU(`��" ���1��
y��hyc�
/�:�9��'o c�RQ}�B��b�p�!�U� <#^ �K%�H���R����r���E�)d����Z��r�����0m-�L��c�r�����\�c]p�ٌ1WRĕ>����2� f���q���S���I�m
�[Vs�!�B(Gxɏ���%c)N�?�G�6��'L�V� � �/��ѿ��_.��j����tSN�bc�-����sMN(���I� �@����R�2M�µ��6��#��S��c��cAjkR8��^;<���T�K�&\יz�4+�@���Y��ʡ�^�m{]v������ݿ�M��%o�_��Vc�1_±�h�J�\��B�sG>��Y1���ϲ+���n�4j�����C,P�g����*�f9z�E�QC�PK*�9*	)u�ھG�,|�D��,�=ŗ����yP��c�
�
@ N�p6�>y�/�]�B��%�L�!��G��c�*��s�|7���W�i�Mv>����� b�0�Y�{dx�f��͏�7���'S	+��nA���S�`P�^q=ӽ�#]��\V�fU}�&��;�M�[U�/	Ǝ��+�Ո�z|��M���3!�ک� �(��p ڿ�I6��K%/����"��c�bxyD;�W�;�_y���L�jl2Ƀ|��	��M�*��9���K��Bv�Ϥ$�e����)�#�#IޣF�G2Z��#��� V�72����"�BL���������|:@��(�n+~4�W�i��Ro7�@O��X��jR�o�/�!���Ruy[���"��B"+4'�����R<;ӗ�B�kU��f�?�ݔì���=�M(?5�ͥ�˭BZ�9���Y���0rP�sJ�̋���g�6{ύ��b��֕�������a���
����+�����g`3<M�&�\�GK�׾~�~�G�����#�1��Ś4��헭1/�=�t���\������B���fp���xvۋ˽��^�����I]�(�&�RD�g��a��i��a�8fN(*�ׅ�`�3�_��U����"��#*�d��ʰ73wӺ�-��vK~L�J��J���wwzPe0Iεi�GY���lG��y�R7�*�wT#Z�'�GBZ��=��\�	*Tr/��_"}���y�LiW����j܇��%�Dg�[��b��735�^*�NѻT:_]`�=L��O$u9�K@
gA�&^�'�*�T8ҿ��fo�:�e���kUW�1���uR�hk���/C�(��>��/pa�]�,��s7'�I���b���h��O�;#����c&�.�����皅�#|�^Nda[VP�Y���HT��5�C��J�r���Ä�����y��M%1Œ��������u��@2�oS�R���-{���SPI႒��D��&W;S��KI$���1;�a�?$�ˤ��,��j�+�k����),ߠ�R�,�s
PɆL�<a�~�k\
��]���m6m�0}jb)A�-%���-1@�?��;v���<�&�#��۩P�Y�t���f�!P�~���ۣ~�ضp��?̇.��wqԢJX-��9�f��ҩWua��R�k]���.z�:_�ݹ����^n�����;_"Q��0����B���5�e,�����5僩n#��1߸p@&�����Y5�ߞ��񯠻��w��U�ٹt_n,���r��h� �yZ#�^��D�ʆ!|J��KPK���CHl��+�L����*���!��I�x���O"�ql���M�h�ݎ�Z���m�$C�\V=�N��`�E�6E��8�jh�U��Ƣٙ�>��Tqf8���ǔ:��%��W�4���{,�O��w�V�o��ݼ���nZe�i�y��ER�!g�6�[@�/wlA�8t�2�S��
U��yg�:���h^b�םj0[��?\;e������!9]娤�0�s���[�zF�Y�oK���Z��h6QU멉a{Fcݔ�H��A�as%��@�H�}bJ�{��*[i���)+���w$�C���&N��Q���߭���(v_e|	hg*�Z���_(�\�Pr0�&<��gN��KE������c�> ��Ԯ��f����[�t1 �嶄��ّ�Q[e��oc�8Lf��(�4��[e7@�bL��c�j����j%@�4��P�v�����I��'�z�'(U�13:,���&�ԛ"��'_j2��W3
&��+m�!�Q �Vt�E�AAU�J��_�[k�yQ$PNg��}E�~�I����;0���=	Ӣ���ao^-�����M	�� ��L�^��(��4���R�u�aK��4�����H����x��?\���)%�j�18�Z��#'��;�4��p����aA�9)$���gj` 1&�H��0 (���R<n;�,l���ln�����/��h����0&��1'9WG��V��\�mGw��A�n-�������,�p�'���)��-Ӛ���+��SjNj�g���5�SD��Qy�?�����" m=��S�f���.J�%+J~��ѬL�M�dC�P�h�����x.	�!��M���[�j!;��N�IY�~{'�&e~w-�j�18��É����}_ב��_1�H��`ҙ�3��lu�3�|�
k顭'B�� oOCJ2��U%m#1I���kz���.�]�&�[-�z�7���')�a�3c��s�9XmLϨv��Q�M#'�M8�9�R0�)$�%�"l�|�؞���#~|���C+�e	�In"�}`毭/�TqAw��'����&x_���q�[fl�J��Rks�V(��6�kS�^BFP$��$άٿH�|��P�ѣ��&������@e��5��Ƙ@���B }����� Y���$�.bs �I�l�M!���3�p�*~��a��n�4([�B_E
�y�b��y6�r�7D��i3�p���-p.�0"py����j�`��<8�\�SYU�����	�u�ӯ�&��oEY�-?3�jk7�b(I�aWV�#�j39Hdϥ9���{�m�Q�XcTu|����S�d�¯p���':��]e�~<�hy���M��S#�)��S2�Ln��@p��A�jzo�δ��X�vG���v�����[��߈���%b��HO�W:ؿ��PC܏-��<x��d	�f���p��@SV�Ǧ�_@ˉ^��ɘk�#`9������d�ê�N�d�C��/�c`��6)�gD`au[1_,Tc	X�7m~�0�\�.*e
uȌ���F���:����)���n]a�|;�)d䗇D �+XW7Ϟn��g:��K�Q��ͺ�`i�f�l+7u�D�'k��2���(�`Rk =G�c��oY�ͧG����0����GR�H�B<�Ǩ��(�ԩ :I���5��2~�k�
Gc��/uʞ�x�鷻�b)��V8��j�?� ��#���/#o1��]R~M����u����eC%��`���f:�7B&�3 D:� ,�bf[e)�9���3�tR�O!eDBp�ާ���'�㿁��1����=IE晰�d՗*�A�v@�HU��?��P�9���
�5s(�� ���[j���H n{��,8�}��!��vy%&/ۑ��>��w����/'��g#7�k�(bE:	�\��$p^mc)µa)�2  H3���)��w���l2o�u���+�A�04O@k����N���ƑTܾ���Nvc0�|���Նq��3��i�dX��D�����Ȝ?N3̡�����˜Ǵ��G�Ud���8M҃���p�H�E�ŕ=+n��6���4\N�[$<��P���4�t�y�)%,
N���F��d�_��0��h��4X,ز���B��mtL%ՙ��09�;/���K^*�0@%�u����p&�{���y������z3%@pF�w��������A�;����q��
8,�t�I�Iby�P�5�/�r�cV�_cM��co�����(dя'<��`�+M`������l?���6�4��
�N\�����]��=�`���2���d��d+�:,�xff�D��XRu�t������T����2RްƉt�M
��Z�{IH����3�D��i�����$A���|T���+������VG��D�My۪׮P�+|6��=`WrdL"11� <�৹GS��jT��p��ugQ`�o␡L��>c>���o��?g,2\auT�=_ip	`r��3���[�lU4�O݉��ŏ��y���w�%w0��/���lk<�p���d�#Zb9�[��s��\���o:���,B�C��]4J>`�IUm��Y�?�_;FZ��r"`���1Sl�  ��#�y��R�3�ö�g���ͥ7@p�h�Tcga�rÞm|֎��Ez�N�W*�{�:���`�a�W�7-���j|��T�\sn���^؜턗�[{��$��{����5S�|,g��/,q�G��;0#Z�]�ԁ2wm�Ko���o���9�4	�yV���� ��z0+@0��,6T)� ��:���'1�!�!?~6�yMkLKp�au�l��L��}�"�0T��~��"�bl5B)����u�L-��=�]Fw�X�*5:Z�����u��|#��1Q�H=~z �vD�2���G�� ��T�t��9�w���R ���G��y������E�Kv��"�����u��b�w�J�:�$m�*�&0�^bPN�9�iRU��ױ���W�iv�a;sq�˶�{���dGP�\^�j��C�3�M�عi�?yxW�$����õ��o\Н���1�;@L�iC���D;��{�I�§w��^tF���1�5{���R��C�;L7����Hk����y$�Ѓ+�{��<q 9A��B�0X���i/�w�ovK�s�(�g���bt��״����̢����"{k��>lI��-@9Enշ�ic�R���������jSQS!��R�u�r_4��/z͎JYe�S�6g�C�&�i�w|aʇ���Š��&��Ozڎ:IS��휯cF�:B�����&^e�� �v�$��%K�<����{P��+�eG������^Q�)M���gO��2�y��c]r�R�N�0�-�T�XlO�
��b�������	R��*j�L���Dv�Y:��Y�8��,����za�d;��@乄v�1	 =����]��zۦ!�-�	?�+G��9�u�5��5;�?�q��#}�̜6�53Rԓ�N���[��`�o~��%\Y���Tr|3a;EV$w���U�/֦��a������6��7��-ꇾ)XV�l���46��4��{;ȴD��ɕ��z*��.KPT���S�����x����<�qR��.n��`�`]���a0�2�,@+��{y_ٕ��C=>	��Ez�L�
-&�@_��]��3t
nfe�U��Q��_���4Ѝ���;8?͕u���T��m�`7��$��>�P\qR�*V�ї�����ãdky��3�Sn��s�o��Ya�q�+�$�)/���I�|���hSj���ϥ=Kd櫨��g��e�|������E��}{Ђ�֝�zف	ԝ%e�Wo�!Rb�A�Y��.���)�����LDE�ڭ��[�{0��&�HX�����]^2ݮȍC`��Ԛ���G�x'��z�I��Tg�V,j��*O�[)��iU7�U'���!�S��>5�+�Y�t��.'�Ǩ`�W�V�KL���J�Z�N6w���ȳ6�X�9�L'I�`�4�5�i�%�E99J�`�Ʒ�,b4tM&��2Y^m��k����{��3����=�(�T�V{��s½�����'7�y�������h3�r�^)>+�;�\r�#���9�@���rů�}{�u��fL�Ƶ�
&�8E�ȪL.&{?�A%�\�{��M�'�� �pʫ���'�E�y�¶0m`6\�[�]��v�������-�=�hG�֮CYF5sY��p
��,�I�����9�T�����N=7�?{S�~e�����B֩Dpl(�U��"��!��P�9l�R�}���H���ke�����s�!�"A��n=���x{چ��S��r�'���~2G�q��l�Pz˘����O�m�1�sXڸ�=y�B3w��@5d<���	���D͑��[�O�RH�xb��⤹z<�=������yBK���wc��G��Z�4�%���sN�e�p��;��u�4�]�Ə���<�2N8z�o��<�P�Qx�B6ڳj/4����V�B����+�����XX��i�Wa����S�iQQ�w��j�B*�m)�~�����J�^�]��#��	/d
/�R��!<��T<f�zS�cZ,<��G�25��$����)~M����_�p�'I�V��I�:�"������N�k�P�J�rߏڹ���3�	���L�qA�R���q��D>�CI���r�Q�:�+�#��8��u��H��?���*΁j��K�.:&L�a��'ь�A9��1l /�Xݥ �����ˀȸ�M�����>��l�C���B?����@�5	�4'.�;מ��U�tA���iZ�k���Q�!�m���9��`at�;��:�����j;����D�S��p��I�8t�%�3ڏJi��'�F�{�L5��^��Ab�W�j^���3j���7M�M,˷f�ЇԪo�G��h�e�eж�B��]o]�X���\gœ"L�!@ܭ�"V��p�
Au���4�0i��Z0����J�x��dj9����[3�L(èR���q�去�y�67�+���:���ii��>Ib����˾7q���Y����c�Ubi��p(�Q	>[D���cnKo�%b�4:N���ƞQ���砛�<�G�������:iM�i]�[~�U��@LY��L��Y�*�����-vv & ��6����,��J1+/�; �3��!|{�ZF�����.��������kr�5��u�.�E��ϻ
ռ_��%�<�_g�ʼ1F���*�@;����f/8�bWħ�L3& ��d�D���di���c���R�R�� teXS��S�IY,���w������q��CI�n�����L�m}r��-fD�17pz��"-�y6�:7(��uJ�J*uO�;����M��8uئ2D��/�Ĕ��[$󚟾�l%'��y��3@\I��X�wH,��I6�,����ͽ���AF`���f
����G ����O9��N��9����K���J�.4SK�ӧ����N�Ra�MS3���g�+�Z���?��:m�Q�7������\����vZUao=8�y��P�����[���ٯ�Ґc���>r���J
'�z��ʧ\�d��M�A�T,���z�?7��Q&Zj��@Ǎ�#|��ht�r�=C{x �����������i��S24G_H#xY�]�!�'�9G�J<v�+&���/�2-��,�n�*{�>�	>`�/���@%�O��޷ �s�Ll���|�w�V�ﴗ�,UC��r�ݯ����q7+��� ����&'�9z�L�Ŧs��9��#G�����׮B��dv�Ht��!-;i'�r}��xK�~?v��><��܎������t7r�l�^������g/��@�vXc톤f}��p23�4Ĕ��̕���I�`0��	�RM��	�~�����\Y��J����|k��39��@�{u�Uj>Ҡ60��+�G U�]���@��>�Gʿ�tP���i��r.�I1���n��� �t~�Z��A5t���"�;�E������^X,+4D���gSU�̚��#(}�4=Hr(�����`��_��;!^�`�Gϱy�{n�I�u9$f��^n�PA�m^?p�=
�!������Vǫ��jt�e�IB����|�0����~B@i�)�a����+t�9̲"y�}C�҇�ں��lv�G�Q�i;�+�ب��\��l�f$�h��M�ĕ�Ѯ�ej��4�<1�G�UHM���$Ga����+��������Z׉�|��\��(��F�E�=_��BO��������0�>Q��|&�A)���?�cBv���bLQ�C<�����D�N�&�vE���6�𙩁��y�'\ ���RY\�}�|&��{�P�W��> �2-G��1��ҹ΃=4(t6���q�O�ķ]�:�v���2A6P��ٻ�^ݬ��E<�*���u�GպR[�[y`��\U�A����b����f� ��oS�
��}�5�/UU��V��`H$�fr/Z&Ua��4R�l�H3�g0���;`7��{;m�B� ��ߘN� g�{jr�Z��UQo�XP����H��y���<�6}v)�P�W9|��Ĕ;7�Ym]���#:�`�H�*���!| Fח(!��ga�Ŷasq�e��ib"���+]�t��9R���t�m`x�yג�����͠���e{���Zv�^eD�i�y���ø(?�-�">r7��lY�����Z�F��|����ݴ��#�g8���_���� ���6��v͜��R��sk�2iK@B �ʃ���U�ͦJ���[u'�>�K ۶3|]|nWS��M�ȳo�U@��w	��"�e�41�NV=}�C�%R�-:���h��uH� M�^|�"�o�A�p|=��P����동��0͵�4d�E���C��Of��,�F-
"e�j��C�R��`^߆�`��~��sP���h����a#Z �WJ�đ��`�Di��1�y� ���r�5����0������:�d�}�A8zT�$��N�E	O`����L�Cfg���t�Z���u��-xoi������_#�aSeP%<���1(l�����u�5qt�F��,lv���Lciwy�)~����֠!ߧ~8�r�Oz����=G��52`���O���ÿ�B�V4<G�^r}M� C��ua^� w���!T��
8�jQ��	��!&Τ(�B�dů��=���63琓P2B��>�Ho2ma.1���%e"!��
9f�}��A���Vf�Y� ZN�'m��A:����z��q]?���O�+��ۋc�h�p �y�~V���Y��;	t�C�q�h����G���׆���?~��w�]!�I�&�T\GV̝��1��H)�{(�S�[z��I�$��pQ��.gJ��т���7���q\t�(@b UА�	�����i����� �G��8���)�ox��>��G���Ytn��7���}ٹ�a�1�K��게�8#��GѵSB�3>P�����~Ȩ ��n�ųS�Hŋ�#�tF8H�4��ĵVk\��=�n*i�%}B��;��)KZ����t���:#(��|H������Y��2���9ݜ�n�1���ǈ�������Ǔ��YkfR�w<7����ϒ�� j`�O���bY��_���]��a��FLcb�y�j�KX�>cER��������ƽ%�:e����x�>��5��4��ȐvBcCg�yO~Y�����u��ٰp��Y�����R��
H�DM���H������� �Yu�!���T�>��c
\����O��+��~��'��v:�����;f �l���f���ט��浃��w[��_�pM0�,�����/f�b�I�Q(��;�+&L����Б��p�p]��fS����y<s��Q\S�՝ʤ�]��x^$h�b��S����퉩(�������"��w ݩ� ��8��O��\S�U���H�%Z<��~G*�\_����A�^�7�7�b7���3=��8�G΄έ��7�?����V��֊A���$�%o?ư6LO?2?�IΫ�`��8�Wk���9���2ռ��9�^�RR��o��.��˵&��$�$��Y~B��G�>\3����U�1ҿ�m�Z��%��@��W�T�}��Y�w��U<:"B�����ha�CA3�
�т�E��'�8ESQ�p���G��@g�	0#���{�V>��6���Q���J�� ���$���j/�81��`�� �8���%���[=���G��海w�\r�{�j@��*P�Y���9�5-�a\r��`�N�e�0��|�`�P�)6fπN\~����b���}ш��_���NtG"�(����r��y�n�#��P3�П�_�p7 </�Ӽ	X�(:�L��=�	�?�׽wړ��壤��* ��1�sXx�JM�ޚ[��F{���!�IW�h#�D�����JI�ӡ�����o������Ha�^�Q;�נX�Ӿk�f�7�E�����\���$�:FSj�yܔ�jS���c2��G�^�	�sv�'�d����~8�*'}�����2H���.�����J�t]g���T?0�>�W}7Җı��/2�W'.��:`xx�xp�8�o��,�Q&[x�A�� &�����@T��l
bSZ�@����|�2��99q�Ϧ�2;	jf/����j�$��Eth�ab\�u�j�/�WQ�'��7p���uᬺ�����'q�0��h�" ��>1G�>�C�S�}n�R˳d��g"Ԙ���60Bk�8	�5��?ī<�?iC�m����jAP<��ޙ�����MУp�~��I	��_�|�;����Yor6�V@�H{�ڋ3�Wݧe_Pί�+�"f@GUmo�cw	�B���U�B��H�.M�lȢ|fK�����_Q.�f��7tʾ����fǨ����BbԸ�G��3-e�R|ڹ�0DE�� ~b����(��~� }�N�]%�ML
6~?��r�c���/t��B0�;�<�{F� ��3k���/V\[=�N���lf��z��BB�&xl(I;���/�<�����7��;F�j�O��Di��,�������bUTH��b/��*�Dq��I�82C�l�A`��tJ�V��l��A�K�O�3L��6Wzs&�D	�LOU�
�����1_�'�C0eC�5�P����o�����
)+�Ut<���\![����ݺ�A��) 6�C3CX��z	�4v�~L�$�Lt�	��Yrg��ϱ~���x	d@�!������q�2�4����q?���=~��B��EmN5R%{��1~��b9���wQ�#p=�7TR��ǻ�񾻂�Q�&�W(�3��e�*�Ȕ�J7�j��3�2x�)q��Fp�л�}�b�M��6G�B�KY���A�  � ��2���݄ΈMaZ���ǩ*f�.� ��Z��F��F�A�j���t��� F�4�DOY�-�ls�xH*�A�|�հ66jK��):Bw��s&"}`:��iM����c��|�oq1�]�p�g�#*�S��ݶ/Sӷ]�K5d�{�|'\
9�c��cRO�YL6<�������84���=�����Ş0�������*�4��!�x�Q��EP_+�Y�����>�4k�C�H����k��7T|5	Nzw���P����j�".�^ށ��j@b?�*�T�V��2�Ҷ��~���
v[�BB1�Q�4��P�o$A���w=Y���#wG��ޚ@| <(6�*�t�d���9T��3�7O�8��X�	�7*��4Kw0P4�k�0K^�g�m��E�l�yf2�
P�B��_�v�|n׺��Ya9���,�{����d�/_��#7w��H���n�U�	�l�Q��lg�0� ����U�1�c�b�v%�f�-��b��{?�F�޴lkka/� i��-Q�	1��0^
5My{�SS"� KN�I��ق��ul�(��\��Jc���Ӗ�����s��m@�)����Z7rP��rlb!�"Ar]�<��	T4@��GW��8�hg	3b��|��Q��i/�XE5��fxk�7�Wmz�^E��M�����o�r�sH�z��+� 6�J\B�mK��%��}<���������
"��Yx��U�=u5E@Gb�')Q�q��F`�T^�^Y���	�}�P�I���a��lW�1G8��~��nl>�^(��s�f=�L|օwdbg���o�'�s*�$?$�EpB҇����Q���8ikm�&�>;��m^m�]���:��@�O�z���~P�>���<��C*�lN�4( �m��H�L{�O=Ki�&�wj���d��6�q� �l���iW7��Y����wY��@B �F�g$+�S[������-��eb��Ί�=\�k�ۘ�=�%���I9����v���9qC������AFA�׸_� b������#*���H�������OX�F:��0����".��z�qF�q�)q�6��PWA¿ߎD���j�S��y�/-�a�tM�¹ 6�̚��Y;�J�;�����
?����k㛶����Cc�z^i���s��
�UJt�K2�_���CRV�i��\�W��,�baM7v�Ν6/v�H"}c#jD&t�C��Q��c+��E�6Ct$ �%tG��t���+W��I��,�H:7-�@؈o�s�!{���&��#v��&�}L@����o{��f\���_�(��e'�:�V�`�p�!vy�{?PiIz`@&��I�pG�����3��F��t�7�����Xw���'H�U�o��ee�v����.oh�h��5�7��c�<p����:Tҧ7�	�4�ت	�5Vs�_��>2V �y�C��s�`;,?K�.n������ӭl��<v鏖� �c!���B?�-GP��������e/��Ts�w:Ytf"R ��9bP��^�d�~Ĭ�T��N�U�z�>���J7�%-���)�ĉD��K������=p�HTn�X��c����b���?Q@0Aw<���L�-]f��U�CJRfő�- N��bը���o���EQ94�u�X�}��C�bg�ߝ��=���lGN�B1���D\Lu @���ߝ�h9Gw�jc�Cqd�!�@6V���{LTo��Bw�"�s�(g*?\Mx���s�_��p1t��8�#�:zJ熡Je��Vv�Xrt�UU6K���-9v�΅�Z���uR��JfTy6<�X^6�}2���0��ݮ���͔�^s������B1�:���^��?��z�y	��8�7X��h�:�8�FHy�f|��&���ċz]ZT��N�Rm����[h��|b�BS?��j<���Vi]��%k�mݫ�r�"(k�}�WI�ȡ�-����J�����u3��ٲ� ˈ��,lk�������.H�������2�p�u��&W
|����	�eS�Ks��4R|���qN4���ף��	��VMp6����g�ن%}t�0+IG���gZ7#qb�NEu轨a�KG@*?v�E���&�$JD�i���ꈄ��2��<H:����o����V%�A�b�zn�G���jcs������^K���=���j���L�,Dn,P��i��!���y���<p4�bg��`���)yh�C��� �bpUUӡ��(`[��(�#4I��XX,C��Hj+t�HԀG�'�Z�#=u�e�4!�k�	��B��@�O�s��֚(=��y)�T�o��L�KؙK�i��fIt�i]�oC�l0	�!m}��8��h���Ùc���{�)�ä�=a=v2��(��Pu���dVY�C��M-|QE�x���P��,`�j3y���ܸ�v��=ϭ4f�9Ü�U���K�!��~�J�Ծ��4��<A,���&��`��I5$͞s}Y7��"�wc�8������?
�����B�#�45H�I��0���NL��%X�jt�h�����2v�*ۢK�����S���N��h���Mf����������`��W���h׉�j�E��pG�}�q�ڂ�N��Ř��^M1�@1��Ҭ��_d�@�[���I�V�4�\���B�wg�bz�����Ӕ��׬�'�s��؂B!�I��evP<������:�1X$�����-�B$ ��I_�"@�7��<e���|`W
Q3�E-D�u�u����F�KKҋ�r��f����6��3����*V��C�g��ͻ�d-U7 	Q��8��p,1��2�d�l7n�p�v��ca���&�#�C�2�7��穙�{��}�<6�{��<��@<=ZA��A1-B��]�T�%e������@xo,Q��A�"~�i ���:sA˲&*��4>2΍/g�,p���ЈzVĸ���Eh�v�!5��sנ~��vv��9��Dg܉��	����$o%H��/6�t5Cz�᫦	�k��V �8�3f����� a�>�i�dRʯ��2�����wnnHg�=�H{�y+�N��}Y��mq,��>�']�i�I4����$o-�D�h�6}�Pܐ�QI�cCWw�n $��\�J��/��+���g�D����GU��YΝ��o��V��b�%���_�d����:�x�qxS�N�a�~�y�)�kn/��t��v��0�*O�TՈ\ي5m�0�x�o���쫎����3m7՝�n���:<��?��˾�	1�ZG��=��x�6��BYSFC=��)d=_Y�|�ޥ07�ǣ{����s����G��Z��F����N��Ե��s����LU��8_���?��rp��R��H���� }%��{�8�i�e��A��o���|�پ�'~��A>V��R��;
�^��w]��8�əl�Ltm�B�����K�ʶ�mZSI�. �O��n�	��ys��������\��	/�B!�^�� [�O�H�ݎ����V�RO����8w�Qk*����-�:j�����9�a^���_�]2�����>��޿�����[A�޿|�7�)	1������;=�f^�ј�Ѹh���5~�(u��6��ZD�����r�x���ӭB���R���|���;��t�c��H����O�~q8~��8/���8���B��̖�_�����1T�+��V��"�_�߸�m���>݈�-�d(�c`+�����6B��ڝڴ�k	�S�"�L'U(�_���WJ����~$��l�_�9���Vq��? �kC��%!ߓ�=�h_���C*y����n�j�w5�?A;|�<��$��E�l��g�X�\�eF�wvu���U#��n��lO:�o]l2^�s�TS����jl^�rYb��b��q�iL�M6������A}�"B�0kuU{�~RRGv������|�A���s'��5!Q�64hW�8�LO��n�PT���Z��NN�;��f-��h;e��V�6rP�k�A��p���l�Cf�iޠ{s�_4+�Ff�Л��T5{vWɻ�����{���&�X��8�Bi�U3Iv����V�ĸ��Q_��MJRp����-9*��F;V:w(��I�$[B���/�����n���|cj��*p�Ňa���V�	�η�.V����>B���%VtnLI��j��i�'o'�:%�]�9��j��_�z@?*%Nr��+��� h���q��px��Uu�?9E�I�z�T�D�,`z�����oT�>�nU�sHtk;��̖n ���5W���<܍��sm^	�E�͵��vY ʔ�iW,&�3E9��0�\�T?���̤�`�K�EyO��ISI���#u]\=?۶�:���P�D�nq���0�e�[��5b��x�s����=/���LWN��S�\���kV��~��S�f�{���5DwH9~w�U����!4S��g�gO?:⑼G�Y�ҝ��V���t�º��D�W� ��@D�U#�!?��g���SK���Ty¯���ޑV�λպWe�
G���	L���'A	��_��V���$��a�{Ɵ��dʈn.Ƕ���T��"61�mh��~wI�ͨg#�� ǊR��
��)�?�Jg#4�Y��r�s���aq�6PB}b�]�5L�ؠ}lr �j�L|�0�5 m>?��%�J�B���H�c�s��|�tI�n,��C@GiOU�����n7}|eg��r��~B,i�<����i�\
���IZ-��hEPy�B��^�l����IK�^�����ҩ��Nk��G�_?�� N�����;@�9G
�ŕ�BGl��)��R����f�<m�v	j[6�.�Bl���l3�nnz�Py:���3�p��uf��=L�Zkz벬��1^'�V�B>�	$g'�]��Xl��XȔnk+ݗ_7�ηǲ�%.�E�<�A�_��M[zUn�NA�������*m	��GS�Ѣ�J�#2��``r0�ޅ����f<�E���#���^����u�{"t��|;�X�2�(�83�����Z�aR.������d
��Ť�h0g�����z��5��JQV0��٠�aHmu�_xf�!�ORKD�Jc�:f�)B鼛�<�
��ݔj����>J�.7&ٮ��(��	S���C6���s�9�j\�N��t�(��� �5rآ��J�sml���qqx�V�����wT!>
������P�)�4w�d�c���_�=z�kB�7Ȫ��D���R�`���v��	?dfhҰW/���$B��h`�o���5�ƭ��ۭ}�EY��LJ�=�:�@/��3D&c���� ��E�KoHԴ�Om��ڲ ���&��:�-�sd�W�����.&���+�LY�ݚ{�+e��|A2�ʋx
��1*j�UAE{y\pT���������ҍ�(��Qmf��٬��Iɕ����Cq[�o� 5������`�+��Gaa������Hנ�Pĥ��	�^�r��k�"�Ng�^o�s�:�Q)���xLIvĤ�u��s�F�x��y��'R�J�3a�J5�I�B����U7 +�H�/�?o��y�B�ܐ-q��F��z��8�4o���A2�r���a��z(P��4W��7FQj�(�>�۶I���	_0�&Ϗ��iAZch��?C�")U?F�m=�����V�����ޞȚ�&�����4�*���L'���A��1j�y�n�Ù@�:ҭ�ϔ�	e%��� �7�F�h�J΢7LA��0@e��Z�9��@�yq�^�pɮ��i8��+�V��t&��;���a�V�N���M%�[���&@']���9�'^E����6)��5�bү�gR�,v����Vc?��*\���ύ��09o�)G���ɥ+�m3�&��R�ͼ;�Ur�����-h����!0���Pn��1^X���0i���\0@Y)b��|�����3�)G+�����R���u�;z��h`����M���f����\�eK�1�؊.@��(���������`�yVpHnJ��[��[��uc���"�Z�P|o���i~=��D���]�4'R�`ax<<d�Oh�{�}HWTF`�"���:G�@U��A��a� �i�g��[�t�"��|8�V(���ְϋ̴�O�͏b��9���aKaH�k��-骛���?�eul��>`��8װP��#@-
@����d���'�����옻�r���VL�P?4��U���L��/��-�.�����*���B��8�����4�܍����#8Q�4��L�h���up���R��ͺ�P�w�#��"YE1vD�r��DE&Ls�B����:��E�N?s�bL��ce�<S��uB�!8sp�z'��v����S�2U���7�������,�C�1P�����^�!����&�	QX���7]G���m����UI���q2�U�S;`&3�ڴ��a���_�Q2EC���vے\Nι���sr? r�Mq�K>ܧo��><0���������#$��ۈ��6��'yz�#n,��mCk�4�\�&�y��Z���j#�Jҁ��9�ׅg#1	�O9��ə��k��ɨ��I��^O���
$!�d����t}��|��eiq�Zi��G_��ԩ�O[�o|����u����l��
������8^M�|������&�4S�������)��q�@4�;��5�s��ܿ��r�� �3 :ue��|�`���,��z>|��.��M���4M��kQmx�1���_�ˈ�вX�e"f��*��i-��s>!�DN��nap�)��S�Y�6����̍k��.�z�XV��6V!5�-��dq�0��	-ec+
���'1�XWe�"��"�oo=�[R�а�I4x	{靴|�
�<�b�;�|����2C�r�;�j�wQp|8��h#�L4�"�-D0zz�%���5��)L6�E�����;Tf<�)u2�ȓW����$	<+'���{���GN�3)�����X�,������缶n_-W�>���M��d��x�J���}�qj��o@�O�xT[4D�%bE�х0�l�������ՠP���{�i����5��M�G�*!2�x��� �m)a�T`;�T�[�ZS�@�͘Y��$m�	���\����Բ[�V|���D@�Vp��G�:�眶-/��&z�m�%���t�:U�wI`Kg��r�/��6"�7bR���2Y��c�.����h��R��qgg,蘯#�D�N��\�Z>���qVI���O�q�������*���[h9oo,�3��&g�Fq�W	�H{���5���ӫ����8t.~�ʼ���k�dϰ'�ە.��������'8M)���b���z�ƕ����;]|�%Z$�9/��圹��p�jQ�BL�G33�AF��]�O��cA���bA�=�,�����S��:|��k�X���CoK&r�ɼ�cE��C�;�C���H���^�;� �S�D��b����
�#L�}���ڤ�7�H��N�p��U��Dn���]�$pI�:>�3�o�<�n��WT!
s��K�AI���.p_�G��p��&Q�gva��ADJ
 V����&-%9��X[]�ҙ%������NP ,MG�n=�מ6�C�����}o��Acs���hF�y��n�R�Ϊ���cZؠ��}9p�u�Bv�����p2��v������76g�I��������I��.`�*�ν�,_˲�YΚ=b&ݕ~�!5	��<�@'V:}�0�C/#�(��j �f�,~��+��mq��.c�����/U������ ����e3St5��BXB������,��rU��)��s��X�t����C�������]偣�c�� �U`g;�v���sߴ�Ke�A��Қ�r��z�?��r��Dg���r��2���"�/%Y
�h[�fMm��A�1c6�G��x]�'��>����M�+a���L�y*b���[�Rujz}rn(�����N�I;#Y��H�R�o�q9�i`��,�M��ϕ��>Ndǡ~Z���.jۊ�%��X��1�g���{Pᴙ,t�e�O�=��9��P *ބ2M�+�N熶c�ĺЛ��0��k- ֤�#�� �����=�2Vl38p9�c�[qwZNba0fY��pě��2F�2H���%BxQ���[��"������gjs�@g��+��#�{��>��B�#Ǜn�Y6+��� H�i�K#}�aG�y��HY�FzA�k3<�O�'Z�~Î��{a�`4�QŜ�~ࠛ�U�m�SnG�q�ƹ
p�B0lh8,��_4}�sfēO�����Q
��8?�z�) E��J\C��w	M(���1(�H������Ǎ���J|w�q�H�#��|N��"T�ѕ0c��*�#A@�3�&N/8uΉ 9l���������j�؃������ѿ�{sj���؀������=7�P�K@��T_������ܗ�Jhy��H��[(�l�	� w�k��T� & ��T�Y̦6t���� ���DC�m����㍾����d@����+�}��w�.���a�w�Sjp�ּͅ3֤dX,F2���~��L��[�0�ZA��@א�㻾CN���9*.�X�#py}s���p��0��cN��<M8�WV�5w^�d_�{q(���7'��+ɵczj6x+xh �B�Nk@:�Co~�w��E7�朵��'z.S��%�79E��'��<�g���
{ې.�B�g������k�w�җ�hEi��R�:S�&0�L������U�b1{+��|q(�Yi��`��h�Ϗ��b�C.��x��O��l�1.�[UF�����F�O�r���9��^��W�[w�Ș�f=,�M`�o>�dߢ`6�>�k�j�b\���O3���=�;B�Wjd�# �Ѽ��+��Q��@�JΣ�.1�+�GSZدV�磖�T>!"��P���x�:9W(�`r�e�vK��K�6eՔ�o[q�;R��*X��/N÷�D�+��ť����_�-�m������_,ajj�Tpj9��Y7�4]�,��}� D8[h��?dty�D�m���׶Վ��c�.�����0�__)��&�Z�s��:V$o:ډ	��	Ў�J��mC�Ɵ�����Wn9��Nt�)1�`�H@WޖMMգ7����*gH8Y��6���*��k3�fk�S�E��8�
��'��2*����N�?�,B���>ۓf3����`�B��H��6�P���z�����W@�*\����aC��?���I������"j<u��x7�c���MILĔM�pp6$h����&e��Y~A��Gn;��*���pV3<:�1=�O�Δ���\s�Nݳ����������O-���L�8��*�S�ktak�7�l����-k{˚���@Ů3e���A/�.�$|5��S�����\��[� �����F3 �z�z����;�K�nK�3��jD�R
e^j�k�\�I+I<~SwM�Jo��DCC3�r�bć�b�ݧ{jc��<t��P:����K(���`��=		{<�_�dC���b��M9�:��A䷭�Q��J/�{JA�W��Ѓ���1�l�lV��?|{H� �}����!z�'ų`��P��-�jy�H�K:���Giՙ���y��x�H�����鞇&h.�Z�2����{Ӆ5��.�v�uY `�4rusſrf���YL?a��d�	V����7�G�lP�	Io�c�S<g�{���&��&�
���Y�Z��Oqֱ	Cpq�M�'@Pc�Wj]r?!8�f�7�-����g�ڢ���Ju�@�F��^X9?Y��{���9L�Fҁ���c?�	�^m�-%i�?�,z����#~#q� z�wc7�)<�|�?U�3T�V�=N�oU���*1�e���&�5n�l 7���:�#Si�t ��NOv�ƽ�o�g�[N�Պ�c��q��x�:u�?m��,��6
�HбW�A�Py��?�ըv���d�-�?I����G�3�P�.[>##1U�sVa���F���(�4���]���"({x����i��`���� �(�ɂ;����$��}����6 ��������v��+����Y�u�+�#Fi�Q���t�R3�lG�:�%S��:�j�뛣�F�qo���rO����"W�\4�������=��q��E��j{�ϟ���$��pP\�F��f��}�7�OƷI̔ຈ��x������=��<M8����c�Y�vY�+4��K<�>K(	�-�<sx5��©�e�@OD6�Cj���F����'�D�a�舒�ukD9�m�0ES,#P'7\���U| ����7�!�YS"�0���iao�]���Յ��OJ�����ei�S��9�����̩�#�
�2r(��p�4[���I��&��t��$yFjv:��e��z��"�_T /�%uՁ���D r������>�q��c�*���n̎���"i��cI��ÄQ� a��5���:���!�)f�	�q��1$p��<�cס#�|[����:I����L��O��I��r���b!{v�?XJ�L��1�v\�#IKjZ��[Ի�9V�U��/��o1o�c�WA&�4��y��5��7�i�3�Z�J{�z���HŒ^4��t �}�8��;���W�*��}�<���{LO��*{_wj�̐VV��cj~��]hM��\8��+�׫4I?b~���boo���dj$��7?!6g�T�N]6ڬ���p+�syd�<&̊]CD� �X_d����_\t��&��x&P���R��ų͎�Org�m���H�c,���k|�O�$2�@��R)���Zٵ��Z
NZ�p A�}9g���0n� �Y��Nڳ!P����5�coJ�
|��r6aWIG6/=����r�<�/#��t���K��>��#��+�8�`E�AWeiҹ���H8�,k� T���j�<2��O�0F�3��|��S[���,A��S��S�pL�
���xO=��W�md: c��4��}(3O��m�̰'�Y +����H	�Dl��\	������@g鿊F,g��3����������G���װ��Iˡԝ�[z5���bʺ*[����-�b�\}��֒��z
m��
q���C���2A�>[?�-�rXDѭ,Ш/���O���i��*@��v���͚��G��Qį&�E�X*o܃+a�D#�!{ ^F۫ٿ��f���=���:kG���KSdѐ������^_i��K9���/)�B��Y�:݄�1yC��ٞK���L��=��1S�:��FC(�'W�T=��i�iha*oh��9���H���5��I;صb��Z�9Bp�(���V�x�VZ
t۵VFtv���(��K�:��
�P�Kj�j�F���9txZM�d߭�Z�S�k���
��*��K^d��DT�����s������w_������l��>�7^�C  ��9�Ć��i��m1�{�M�:�g���DdCR�^gS	&���8����^�t6p_�m�[��<��|^����x:���0#�H�#���>ŋ����)��.
�0��E�77"�g�X��5���B��@�z�_���9�[�����}��^`�0ix�L��F�#��y!�px49쇎��*1��(^����ﯬ�ۑ!�������4�f�0o���b �����Gη7�g���/M����#0������$@t7�R>��6�Z�9�Ng�>e�3��P�[L��E,L��`˪4|α6�vT�}A\a_�#@@W�������s]WK
m6���un�+�|�r��.�Ԇf�NWȧQXG�|��9���G/p��M��Ҩ��S���m�P��ߤbf���D������6����r�/1�b$�ڰ�2�#����Pk�/y�:��XB���99��ũ��,L�D��ǵ��5����̱�+
7�� �}�k�7~���l�h�:^.W�b!�
����+���}F����W��l$T��zVň]�J䇅��ؙs�T� �ک@Ɍ1�A`w�M�����O�t~�U�c�O���a~|W�W�j�i����2Iaٳ�.��߳r�p/�X3�R�K�Yak�6)DkY{\m;�n/�S��Ns�Ņ�>�4�C���y���`jWr�c6k<{��@W�{ ��>aH�P�>�]��}���)��"�X���m��;��HI��}�`4�y���c�����Zô3�`ohɑp��K�y�E�C�n�
�0�;��Й��� 6���F"wڠ���Ǵ�W�Q�oҧ"[�W	C��+%�PeD�����T�G�:�r�����1����}��J�k��赜�En�`���:�k �e��yC=ॳ5�*����Jb�	v�#��J�Oz'��c���f3��7^�dX��R���W҉����֞Z���:@���4��ݷC�[�qDfx|mE1�{��BnZ��W��6�W�8O�㜻�Cs ����8V��i#�/�B6Z�Q �M��Ћ�<ϐ��o��O'G�2j�B4�D�?�+zY�!Q 
�������`K�Ɖ���&�& U�����"�)2��oSfR�T�|�N��+�[ΖW����w-�ޓJ�`�:|�ඳ���>'P�Cq�nf5S��@���7LF+��5����/v�����ip�ۋS�[�w��|�D�e������j�;T�3eVg�2E����7v��ӊ�����l��򯉶n�{��w�4!u����-�e�k��(���pu0#3)1	.ﺶH�ѷEd/U&�/~-�Ą��!
�T�V�"�]/'���21u���sY3��)��Kh���ˏ����VV+l�Oޙe�ø)��QB '^D������` ���qt Q-������P��@͒�T+w�t$I���.���M��Xܑ�w�H�-:�AEi��K��L��?n���@Gqk��[�?l�3v)N��.�rUd��5�����-]+Y:��	��.�si%��3[�S�Eic½�E��<�h��f�ӒG�QD�EK5�	SxCI5���W�X_{�G�J�͉=�w�QVC��z�?Z�щ=��JM����IPĿ�yX ��g���(�L[��.���ݳF:k0ߙ�~�=](��l��^���HH�V��t�c�φ��|2~� �k��~���s;�-̈́��ڙ�S"�s�~�c1^ ����p��Vg���w���4m�D�#gF=�d_�(�_P��fh6�J�`��c	�w{��X	����@B�f�F�e���<
��\(Q��Ja�����Z��>�@^��@�1��K��o7+0P<G�o/�Ll7����Yv�J�����l��P��s���~�$<��/��s�Q]~���BQ
�!qŉV��'�宖S���	�$��M��=�z�z���
�n�o<`��������k��SS�>��,؈��1;.�����g
1��"O���W�D���su?���>�4K����u�9nI2X���`buޞyu�v �͑{X��d�]����to�ퟀ������^�2W�}\�ˬ��0�UX��I��<��kM~��'�(�i����e�2��!�"�,mH�H~�dwUIT��)�@4�͹�~�[�]}S2�6��8/�"j�ws(Q{�����`G�G�Xվ.u��_hQh.�����5za�l[2=r���
A���=/)zC3�%s,Wa�Um�����}�t���0@�~��[7z�ϓӖqDf	eJk�qi	��!�y|LW�콤6��w�wI���WǏ-0�:ڦ?%�=�1�^bC��Q}`@x8�m
y'�i_:�щ'��e���J���q�������5��'X��+�Μ�.Gk��sS⥪��ɤ��5KD+�j�=pa~���ta�Lm����Dag}�q�u�Je_�J^�m�9���]N[C���\GYk᷐[R
�l>�?����-�q�B�$��dY��� ����"�Q5�:���S�!!��úҊ]�����W'Psf�ּuά�Q��u�0(�6��Z���F,h��ŏ�t����BR��N��!�s]m	�Krk�}Uò����m��P�tf_d���_zV��|D�4�(���1�wR���F�+m��XOڜ/Ќ7�/��ek���5 �����bڗ||��;&�Z,������@O�</�fBR�8��q���(.���6��6@��M3�Cp��mi����=�J� ���G����:ڙ?ꪥ�9	,ݗ�����I�l���&�b�Z�8��\`P�B���)��Y�K�'�Sw+��+ɍ��ds_/7�a��`#v���Y��Ly�*����u�ד�E��+{4��oG37��ux�� �������_[d�5w�P��ks[K_M��3�)��g�Y�R�^D쫱��eA�yw�6�zy���z�k��x�e%�.����R<m�) �����Q���v;�OTNO#��o�O��b�w�Q<>T;�OӢ�4�Q���!�41�	-1�5M�	��P�x.^�Z<�1�:=j �܆A��2�e����u���ύ�.�1��]�rN�~���>���;��4˕��Oj`�����I�z���*�yx]jfܡLK���6�H�P>��䎻���J;����ߡ%���m.�)�~�C�_A��_x�a�Ab,���D��h�"�Bw�ޑ?�O>�?��Y�2r��LOz�c��` ��:E�k�h�y X`U�mn�>�CqCs�:
F?ν� �]��W*FLG����ڴ�_w⎟�3��&K�۽k~��RԸ�>�/֛�\�����0W��ٿ��_�*��o��M����r���p�q�mm�~�t���2]EWFq�O�?������>�&I�h3��D��Ǭ�Q����b���+�mS_ D�ô(���1s�|����G��O����`�AM��;��w����2	�i�=��R'e�Bm��L�����FF��(���V�J-B���pe�+%�+"�l����Ȩ��i��i;J t�1J�1|���Z��/E���z�T^�K��ա�ݹ�mxK��΄��' ��)1��2'O�ub��o��W�[�������%��lCE�ƺm��N+P�a��센?@�r���������jX^�
�y^Dw����Vs�$UV�: �UCK�8��N�>;���Tp���@p%����t�k�	(�{#�?��ME�����{�'�;�C��|��"X�1 ���M����������)�=j�䱘)a�׃�
���v��Wd2�p�]p����er�P,�5�-��>/���b���ࢣs{��'�"L`�YO�`0���\Z`ZY����GD���W���2��*��>9�i�_��%�*��@��Sc'TW�/��(O�<�}r�܇�#X�k׶���lV�_#��W_ܗf,~y,zG$x�$|���:߭��5�6Vu�M�z�|���OPeV�8��e��0D�y��-uy!��&KBo� �溂���`b�k��>��&�BE8T	-_�ݫK�<fK���7H�S�����ս�y;�7``U�z�lhѢ��oBA}�CX�"
k�
�̻��)���1�3n*5�	%�e�_�wvJu���[Д�c^7�0cDq�摱N��l������C��W�ٙ&X�C'͵�����xh\S#�S��G&ur���j��(�ׅ�C	�M��n�����@˗'�+�`b��]RfI��ɡ����(�����2/V�v܇Y��A~g�x�
ҋ�%��-K ��/�ƅ�h�Ɋd��y��ב�)d5�e�{C����}��+~P��n5�CDb�s�ܦ0&��c˾_!��񄦜8�`���A��`Ab�aS��ףg���&܃�|���лB�ps���� {:E�430@$ΛfOwƧ��N�3"��^T�+�Zs]Y�i�j�^q�x?��~1���~j����ϋX{%^�&�]�&��d��$)>��8XV8=�1��pA����6��;yM!�7�!z|��o&m�}ݛ_�ɠ�������rD���Q�Ag�ǶI0�\�n�0[3"J�-Df��E�'��*m�y��ϩ�H�9\W"FB�J>�G��+k�j����B�5[�m�ޡ=����4\�)�Q�%�N�	�l$PJ����^1ڔ<Oݩ�J���_@�lv�g��U\�!���W�ޅm%<������zDX��2��'�sc�H�����͈�\��Z&a���A�2�p o�~h��|R��v�b�NBr!�^�Wq�:�Q]7��?1�:s\��w)@�
����`��0��D>S�� N�I�	�:�d���K�}�Nv
E�3�Ƒ���l�O����Ā���
H[؎�X���y�|����R="ѡnwX'�:,z 3"��`�5[JaM%b<Q�LB�����
�"S�I�S����Z'�p)SJ6���&��־�wy�8N���*��!i�W$��RacD�I�0��}���E��d?zu�ie�G��\�B�`��O?0]_��'@5���#�Sp:D������V:%;������_���A��N�{[�Ŷ��e�ݖ�w��q^��&�Õ����Ŀb� ��O�뾃����ݽS��q��q��W�1ͬ�_46�`C�׾!��d3��o���fg�k�e����2�G���7���
RVpP�F�O�^��2��-J�:�Z��#A�h{�[|�"閅��FhZ�����5�ʈS�0b������U9t�s��d����nr��s�3�]�����3�8��L���,<J�E*��m���G҆oxz�*߉r���~kr�'v
�D��a���G^1�f��](�����h��s���pkBѯ�J�g��rOl�^ތUSK���@  GL&�/�5��8jd�V���w�l�;�-��.cU��伜��MA��kA�+s��� 5��Vӫ}���ȒU�Sdt�HN������9����^m�J�Y��x~��(�*��o�V�����I�
w�����=C�H=g+��O�+��1I��h�9I��,@<lP̕�%��g�H��W�uѼ3�y{ ��Q�h��I��j�%
AZ���dʹ��� $7{k�H!�z$�|�0{�O`��e������R:������$�x1Q��NG
��2�s�@�	����J��r؈!EF�w��G��o?�s��4���.�R�ݭE��g͉ߣ��-ҁ[[FQ��u!H;BK�����SUm.6�D�	�A�&ئ��(�Ûyf��S�(����eP(]K�������٤��#�M��.������t����/'���`��ϕ
���
>����3'�����)- ۹�<�|���) ��֒��:�Q�"m����eC�����C;��ؒ��0ɜ��Ͽ1���aL=��>���/6�``��O��c�HF���,����ު�b��
F���� ���6@�0�cE0��g���D�Y��XC:u�����wGx���.Y�b�*b��y� sJ�Ci
�ӭ�)�=SP���ŪD�`��~4LY�@G��|�+��WI��������+����U�J �m�O��x�a�Օ��TI��s�d���J�i��#���Iu�q�W'.�)��B3}Z�o��H���p�n'u�;LT�������%�#�`CpJ�Xdm�qSp4��W�a�3s�	Tl>9��vꉌ��v(l�j�k� �	x�X�<DN3�ř6�ug ���H��(軱h�A�ƎJ�xI������/�_���7#E�l%_�Z{��m�׹�<�Gź�,1q����+���^h��b�Q遀߃ϛ�jV�!'�0��U�}2����e �r��o^�/�=rhuw�pҜ`n����C]6�a��.Ok3�h�;�MC�^rTtsy�Ԋ�6�S)�)`�ڹ�Q�$�3��=���e�pe�s��J!F@��~Y��rU���@�'��6���)��آ�s� �~�,��ޥ��4������^%`ie�U�I��s=��Y^�[*�v�2&�1Mq�R��D��$����z�
w�S�X��ik�>���&-|�A����	�S�ܧ���$�$��|9�(F��ȍ�4�*�6D��
?լ�m�.U��2�'�3��Υ�a�t��ӕ���$a컻�
>.=�t���8������/��e�7�qs@Q��u_O#�B����Q7��z˸HD�%X����k�M!�sTz��G�\�� ����bI�}�w��F[����������{^��w��ت��[!��JJ�����n�������h8�������`T��l0���`�Ｐꜫ�G�O��H���hA{0�I~�U�����K|�3?�_$'���çª�����
��|���^�;C2���C�DƗ�$礘�*�LLD�j29sē2�v~��T��^ttR���Å�#�yD�K�H�D���Z�y5���#��ӔWGiu{B���r�]�/m7��+�A�bdhZ�㔋2��+SZ�2�!��Q5�Y/�Q�Ҥ� V��\�����a�;��+2���AP���N�HI%@�:����{L�Q���-���0>X�bN��j �������!��x8���4(%�Q�0ac����]��*��?�������REH���Z�g0����EjL��j$1���ψ��Z����J�İ�gvo^:�fL/��p���;�z9��Y���N�Y�z���� N cӛ�.�OB�xor�)yb���x�r�@�>�9�\��]�i�� ��o,���<�5��"��ݨ֮,��&�;�T䡌@����o�'��<z667�v���ZL0P.�O`��!����p3�aqۗ�B-�o��|>ȳ���+�˙z�UJ�>�
���uՐgA��ȕU��ɕ!�v�O1�����Md�2�O�|4pv8��k�G���;���9j_�PW��e��¦���D��ƾo.J��/+��m��(�k�ʭ)�$��/7��A81���_6�5�ۺ�;<��nV�� ���0`�ce>v�Dw�&�r;.�&�����ѻ�j�9Á!��F`�(��C�cyCF+�Q{�rH#��ՙ�t�\�bT���F������'��e� ��Čb3�;���n�r�x�4؟����ѷ�$������q�C���v_������<{��P�A&�1��T�)8�	�~���H�$Pߠ��`��y��8��;F��?ovyl�EvMK���bG����U֚��̀�&��hv�QE�>�0��Ŭ��c؝j�RN�_�$����k?SQ2�,+���?�n�d$�W�W�Mt���K��S�����+����y�YV/ޯ/�{�g�S�i_5��c2�?�dcc�$E��X�Í��\�oa��\`J�=�
�'F��x��{��D��me&�:C���Oq�7�1�O*	����1��"a�b�}|�B���K� ث따�x��e%J�_<S!0g��/�������
o7�����"���/�����B<+tw_����A��-��翧{�x�a�����̮q+�`Q:���%�@*�*�ɏ}{�m �Ori���)|%�n�W|�.X�����[��`�`կt�535{' �͞]r�+�Pe�¶Xl�#��6���D�C�M��d���<����~S����<fۊ�	P'K���J)�Z�ޣM�,����+�E���A��U���l΃�Yw��ˈ�<��TG�[�:��&�
 �%�{H�awu��>�0~�Gȱ���
]��`�m��j"C3�p05�K��#5xbU�v�O�DH�.�|��\}*ZRRj��i�t�Lg��/�7���D6�}���X�ey�SBWN�B8\	�J)Q[m�bUx�ۇ�v�~���p�2?{[Zl2��N����ޜ91�<�@}>5��ǹ,�=���1X@���3��<=yM�7�*'����f��tA�B&o�1�Ω~vw�.��+�[� -�9�+�X�0�_ܞ�,�$:.�E�ֆ\)���mg�k�R�����ۛ���[`3�O�t`�Ϡ�N����a!\f0��4\��
}vSn��f�RO%E�bO^Us����mF|�x7������q�r� 4}��Nn������羆�ڿ���=
D� :�`[H�PH��l$�]% ?�'���lG֮+}K\�G�l�Y�c�'"�m�ۻ�2q!z��B�H	;���o���F"�3$�T0'7q��n����RR�.�ǲA=�eB�wf�hN�;sp ����n��x3Ejd����^�т`=mflE<M�2uX��bŴ��e�1�E��](b�d�p���D�}�/Nܭ�Z-����n[���I��g�7y�z������}�㗢=ԑ35�3�ȱ����we�q�Cpx�ɐm�b��etHQOv�gTH4���$AY��%�lGT�����3̉�A�)��n��o<�>O0=5�~�w!
��E��4�8���s�.w�i�!o��Ň���7�������6e}�K:�p�K�BWCE�}�!#j+#�6�<�%��9��b�e*���c�����V՘�c a���i���ñ�S��5���W��]�݄�MGj=0 G�:n5��g�Yх{y�!.�6�����4 \;,5���{k�6��V�ZVƯ���C8v�ষ�`����A���ߣ��y��ڥ�y�a�O�a���Hkٔ(j%�8Q���9f^wS������[G���������YI��*���N��8��4��SS*BZ!z�� ,�'Ж'�ӫqp�d�<)��H_n�|LO_�l��3�8{nk�c����x�;@I���ָJ�{�7�@�_����T���HFI'�r�ԃa �)����ly�|��(�{0����;[��u�e9ѝ��1$�Y��m�sfĳ��_�:b��6dH��,��_mX���[��@kI`��%�~gݕa��{���J�/��� �k��kG�v҈���B�2�c@@�Z���kJc	\��$V<����7,v<�IƇN|�6U5���G��
�;����dO�d���>�e�h7´4�����-��d���^��6h��`w^:�Y��u�.���a4fU|��æ�k1���T�ҍ����3�ēsPӦ�\륃tΓ-zu7��!g<�uG,Z=��;�'� _I�YZ>�Bl�F��V8N���5�w�PC��?�m~�M�10ֻb�q���L.�=��_�˴=��(��n�2���"0V��X�+2F�S�y����x�aϭ:�ݗ�!���@������(��Z��H�8[4L#�[��'Sa2�*���"�����-n���n��Y+V걃�w�sb.g=���xA>R�\��C��gV��
�5���z+�� ��8��~�p#V+�a�2�����r��B~�o�Y�*��u��̯��;�=�<
�G�R�b���6<ESTl�ǂ�ɫ���o>@?`(��N���<�<$v'��t%��ڐ:�U�>#ԭ��4�w\�/h��s#k�	����^x8]���׉:� �D��u��梫V�i�\ph�?zf��1��)*.b0�;�@�ƛ��2
a϶���r)���3��[���|\,eBbI�y�//��)n$!��3���U"��3����Z�%�-!i��-���"o�\:��Y#h2ra��/ QO{� Mu����HmtRV��f����	Z�̶�|�=x\�6&_��y��=���8o��LA�6h6�D�=��pn��������Y�1%`�=�{\N��q�B�Y-�����a��C���%S�����e�#o�|��F�v	�-��͇��Kk	W9oI �֐�S�|ͩ��N#���~Z��b��2>^^��%��h�P{ns���5%��?�O��/��ә���*����K��#��}Gs��8�^j�u"n��"Eo�4@#�?JL��m�0}.wU��4�<mr����/^M�}R�Dܵ5^������q9�"���/�"=�ZDbz�F�7Ӳ^W�GCb�L�j����:wL����~ i>1 ��i��ڞ��~C��D{Ɔu�&�P�����_Sa�u�z=�׫�麨�j �J�[.��/E�ʉ�
�odY�-�=�Vj��Ⅰ�h�Q"����1MP[m] k��2�ʝ�^���"���l�؋9{�-�X���� ��OD�[�'�Y���/������*P�Z�=���2���'���C����e�35��L�E��p��z�W�q5���O�X�^������6�j�;o��7��xf�����ڊi�4�"��r�2U�?�=�T�D*��].e�t���J�5���p��r4�HI�ڜ2�2����o��8�}���'���f���#��}�Zq�HNJ�E���R�Y�y&�Ж�b����h	HQ��2>���+;K��U�3�����?�e�%%�L����C8�9>�ܕt���Y�rOw���L��3�JeOⴶ����%6u���B	v&do���,�-�N�]���W�ExR��
��4},�h���Uj3�s˿��jc��O�Y�pV���k��*���X�I K!mr� %��M�5Q��XC��Ƙ[�wخ��0�W/��.����=�M�����,�cu�(	7�e%m�m�����d�n�#'��^���B�a?�#Z���thh�6�w+zBғ�b���1#V�|�W	1{�cxau�iO��q��z%e�����Ί,����*�\xM����
�jY^���f���f���
��kX���6�œ#Mz`�	�T@.(wjr�>��b���&=��Ka�
�Wp')�Q��w�!]�>/
}�V�k���߽Щ,��Rr)�i�\�����$���~)�R��2PR��4a����E�kc�ٔzQn+���������'K��P��2Mr�؎�V��jw�+׶���l��y��R(*v�6R�f�S�%%���78
`{&\q�Wվ>���+:�ro���k��n.�`8J4G!F9v�"
/,y�_����h�q����	0�4�ؑ��/�U�^�Gt�5l�a��{Z?�+�H��/���?+3�'P��w��m��Έ+2d��^"f������X�o��
Rr[�*��g�,?ZY�r��X��]��Љ�M�u���B^16h6��	�hp�|?�)��Cs::�fP��w7�,�o�A��Ɓ�x��Q-��M��P�%�,M_o�~s�kUg�`�g\u�
��ڿ�e{��v���v=K<���B�O��썳�|��3�?�޵#��3�:4|X$�El�Z��/A���ɵBՉO��� >�G?C�I�=�/qz$�>�D#�uڢ������Ȕ��#Ʒ�z�t��f�e�E�ɪ�,��6�@�ߍ=�ካ��>��:�x�?U�7,� ��y�5m-˪A��';�W��r=
m7Y����!��0џ�ζ'&w)�<0DYLGU�!�"��I���a`�{L������N��:?���1��g9PB�v�2�=W��H����irS'a�~�>�|�������	Ѩ�\����//?Tl����'(C$:"\�L�x�����#���55�o^!9<ܲA>��8��)���SH3��#r4h>��$>��/�t����/�Lp�)	��/ER�t9H(Z$��� �*ae�c����T� 	F�%O�M=s�� ���֞#�K�]���	K����b�ix}r�gҼ��/��h��hm�U<�2W�Va�Z��P!t��&©���d\%��U�Vf�7��<�WXj���o�����OɁK�C0'oV��]W���[�u�n&"��c�~�{Ʀ�<�Jy�ʽ����=tĭ#��_���'�f~ZT�&8B��$�#;R�%6V���bרo�F
|݌�]^�r�����.e�V�Qf}ǌ׎�y<��@
��̧ڊRIuBn����V��:��Y��$X�HU���I֖�����k��͐��a�,�C/��;�s��8��� yzs�L��L���uI�^��t�ޕ
YW��8�Ȫ�r�w�z`Y+�~��nm ���p�1a�pdV wOs"�\k�'hH��HQ%{02��15�����Q�2�r)����� A�������z�.M`�)�t�bz�X^a�VYl��]��$�����~��]Aç�S{���@̖���8ڶ��VF^X�>�r�<�\�>�r-�8���ڭ `-�"%�J�[z���ԥ���]p�H�F�W��@I܅j�ݒa���f��k��B�D�uU:eI@��U����O����T��J��t x���xD���oAD���
G�3�J�҇��	�F��!��f:�\�c��+�����X�&(��Hol��l��Rh�8�+�,��sNӤ~֦�N{����7�y Y�)+�+i�~��8��AZ.]�K��(�@��mA�P	�t��~X�������E��oeBT����clzKq̵Y?b����:Ǵ�B���>ˠۋ
��݌�$�����F}��R��[j��)�N��mhI��u�hi��)�	�1kv���DM�ܭ%�r)�V"5�4���H���&��|hڐ�_�"�֎C������8�]�����&�bO36�ŨA�X�*@��{�%�F�GکM�V;5s��t��Ŭǵ`p��*hSe�b���ק�Q��l��v�po<H���>��D`*�B����[�������@<��^��l�_���#��"-��L-�wU��L˪7� D�S�VP%�Vָia��yvW;*��B'��"���%j�q+���ߚ��jQwY'���N��QN&�u��v�D�14,�6G�p���NogF}�����+�_�ɱ�)+��
�b�j���|?]ĵ
�x~"�0��u�l\w�����uj�=��r����z�rE�����G���7��gV�O�83�_b+���i���VԪ����e�G���)pf�����wl���i�#d=��[s�5�Z#(�?w�J'z���9���N� ,)�VGs]|�K6�vwN�ak�a�C<P��Oq�ԌJjas�!)��1y�%�|�f<��ꞵ�o6{-�l!C�Ի�c�)8t��%��G�7D��g�q����8���s�������1MU_��#@�n����O̴H�i]�VԌ���j���,Ũ&m���O�zyu�Z�뗚��a7Ɣ���<2��
񕊰xN��6����Kg�)��\���6_,@��{?!�\�Q�RUO^w�B�Ũ��Z�5�&s���i^���O]�f�WK��Z6~b{N�����=�	�}�;�5�P����0V�Ev�h��`EիwT'5�~�_2/c��4M5����|��P����l�zt8W/�UˊMy���M�s�C�/���8o��|�ɤ���u>BD�=2���2�%Tʇ�" ��9@�z�Jp�I:*�]PI5�M�m's�FZzbBd8����������?�}�)YH���=�ݹ�J�h/e��
N������~bq{�`P�P��s�fO�{��/�0�l%}���:#G�7�?���㖓��k췂@�4;9w�~?_�l��K~rQ����Y󦋈�5���T.�������Y���:ZP�d�F3T�w>J�Br��u{G�:��E��<ϯT3�����L�D�\r�0�ʬ���Zg����v5��.ݵʄ����L[���l����,�;����f���v��p[,ND9a}��M����̡�DH0}��K�qR^�/jL�{0#�h���*����3!x� Ρ�r_���J=z^�-th�x�J��$9 �`�%��;ĸ9i4%��NX@Һg8�*`��=;E���;�s�
s=����7xʬ�?@K�~Vd��>i�-6��E�K�'�E\'�h�~.�_˷���ɞ�*E���'3﮷� g��÷;q��a����{�T5���G� `B$���f��M	��m� ���	�?�M�7����
�����c@<�(F�$:&���L����~�Y��@7Cù/�,	����������˨�t�eH	~��z)�ک��0�b�G�+��~B�-�DbF�X5x�t$ s~0��ܻ����%��@��?a�B�P�RŴH�e[ʣ�`��<(դh�Ր��k�b��y>%�+)sf��H�j�$��'�+�{���MI��n��)�$+��^�vᄐ�#�?3����M�}�K�L�핱�T�;�
�C|�M���R�43<eu_��צ(�b�L5��< 7I	��0��;�wհ
/���y,����s�ĸ�����`������Q���5n)ߪ\	��H����#f\���%B�Dճ�$P������K��nt|a�����
�<�[<M�cb`��:��h������z�)����1�8L};
F��uI��:�p8a`�l<s���[#�L"�b�~�T M�/�g�c�}��a���J���}{��;��W*�=.�N&�y0�k��ݺYG��YQ�Us������/�,�~�jU�����rه�^V��c[�)�j�;뀓J��L)d�6[���#�]���&�J����[I��g/����I!-��V����/�a�lP���"C'��8p�ÇE*�-�������_����);ȟ(����o��=o|	����ЍX�!lv���gJ�w"XIARW�CWx{����N���,v?������O;dq�Z\����c'i�n��� � ��SXR�EJu�A�e	@JuY�W�;$2aR���L���p�5!�)H��x �x�����)�x0%��4��-J�!�<��Z�\Fz��ls)�Eq�6��]9�t��ԭn�j�����I�G�<�bb$�1�pl�`�j����Ɇ��NE�=k���Fv��V� �]ra/R[�����#��GB���V���a@:F�s�5���}^^.��;�fŁ�j�(�q�� ��vS&�@��wy��Y �c��{��N��i]�8Z�+�:w�Q��!��\�� ��7���*�XE�ykh�/;aFN�2G��dа�]���]L�WSD{����֏�y��'��L�K��Y���eZ	 ����f�Z}I��Ja��{A���ˮBh��u��`�g�ˇ�լ��	�<k���(>�弭dG�ojR1���+���J� �l4�$
T~�̫��VfHxfߥ�v�x��D�.�)���+>������q`��'xI�i�VQe ���#��]�%:'�,
f���"4����ez_P)_�05��Q.i��Ʌ3T}�T���k��k3/��H~h�U��h�6�B��i�͢�~h���"m�y�D�fí��y�P#�%�U��*����NmR�N	�xz!_L:x~�Ӌy�r`V����#�2����l�w��x�H�����8�ę��$H0�'�� ����I ��rvDZ+/&4@9݊��	U6�*"��6��?>z�G���]�A[�� Ä�q]i�ȍ�U�P]5&a�0���c��Y�v����{��v��!��'{�3�M:
��&C�-���4�~[e塞+6�0�Ŏ�|��AJ���SvzTy�3��A9ߏ=�&���"��n�����0���HU�%>��B�X_=7�N�� �}[(;Zk��*���5\T�̚Y���5Zwq�5bZ�J#a�c��LC�߃_��cAAF�od�숊����B;F���L���bv}�����0=��wO����<�	�_\>�1�Н��5��������wI_XD?���K�f��r_�T ���9�جv{�"A�6>�`��!��;t�K��<�7��]Ї ��c�_�M��{̔�[�h4���0�@+#�&����P�v��!�G7�ԯl�4��S���.8�$�y,��4@�9�?դ��ك��,B��F�<t0O����HO����a�u?��Ơ�A=�k	�1>�D,���A���>��u�}��������T�(ghGNn��tTÍ̉s�q)<A��*��l`�ֿ��K��Ia�u7��v{��f-�TN��~��Q��C���K��DL�k!�cW�����'9�!��/[I��b�^l2�&�c ����1�C��3�И�'��HI�5�u��.z��鑓��x\�ӓ�o˒_У}�3J��h؈�,
�t���b&�6���Ʀ�W,Y�mOk��$�=�>���#ˣ���ZG��=ܘ��^�Җ<�6_�F�7eA�!���J0��K�S,Բ
, �Ь���{x�eKڑc4&)� �e���g{"1�L^���%EI'���|����LꁬW�iحœ1�8��5����dߦǈ�̮ʇ�v�^+G��W(�(��\��oXw�߰��9(�t��Is�
�/�[Ô��ȹ��e"�����=��+��4�����['�^���-V�>(d�,N_+�^�ͭ�G[@��1
b<���P�_
t��wkEP�@dx��낮]��>I�y��{T��D�o��}Ǽ��^#n�����ٳ=�MupK R,�Z�0��kћ�Xﶔ ʽ��ۣ|�jzs����d�=��Vθ�^�Y���y���o��o�a�.���7���8U���
�*mͿ�8�tS���
�d�Ȝ��ۄ�r~�÷ruPd�|����Ԝ%�E>kj�D��>4�,������s�������<��	E��@�0ꮡ[u�\�4gCRق�Zc�\�ϻi�ؕ�.uV��O�!��!�F��|`�T�R��ɟ�,Vp��0z��~V.h���c��an*aLAss��4b�����`��V���	��q�����Q�clJ�O{�!G����b�m�jfbH擛��h��q��1t�f]+n"�#�������7�9�D,�T����h�LO8��±T?#TQP{�^�{�;��Pq��ؑ���{���?��*!�-XE7|#6�\��9���9���Z����z1�^ĕwɦ�^��Y��
A�)us{��G���<]�˥~�	�Ӌs�����<�+t:�8m*� HyI?�_�6E��L!AxC�88�l�@��
��Gc<ZI�E�y���]�B ���I�C�g�/�c]��
iH�C�. 9,y��k�Ԥ�D�|�3��6�d�t�Ǉ;� I��+�{�|�Q�z��}?g|�#..#1���K����Զ���*
ٗ�>��Ӷ�ߖ�е�h9���p@��U��M���oЄ< /��N��b�k�y�=�u�ͮ�6�q�����-y�N���9�X�X+���4Ʌ8����6�),��+�q0Fk�(��[ aA�۲�kU��ffV��9@��K��!�|o(���bh�%J��9< ���y". �`� ^&�N��n;T؉ek��n�o��M�J�}>�(����u��u���ƃ�1 s�T�;�G�dؘK��B�\#_\��x ��Cʞ����'������_YB�ȅl�����]��M#�X� oM��˓VᲗ���ҭtK�7/i<|�/D^�����{���^��F��x|�2����*�!��a{h�&L��&2	�"O/m3�n.��2k��@�~~�M��n�;Ż�4V�m�SŜ�5R� �����6�%w�o�b���Gזp�2�ȯ6PeX(hF��U|f���r��l�f��d��t��,knSV���P�mv�̟C�S]!d�C�y���7����F�0		���M �"Y�ʰ($BQ����a�+���Vs�H�
f	�2�s0��kq�i"ݒ'u�i G2�֭�R��(��oY��僌o�%��c�Kt����<p����?�e�:F��l���{�Z������J!���!g��_�c�8�R��%\ڴ�C��s@�w�NRZi̳��ҏ����-�w�^A�6@8��$�������d���}j�N@�婥����0���Y"���&��j���A׌�Q�Z�����o��d��WY�l=UWN�a=F�����d7�Gf��s'�T>�.}_�����{��m�0P�A����
���-��!E�����U�F��P=�ސ�٢f����$���ީK 3�v�\@C����붕#'�j`����~p�a�;<�Ħd�~L
	�
��ef[*� �񔤉��ě�Weg3h���lk�(mX�YH�
d]^�,��n[UQ��m�{�
�F腷gYq<�|��f�}h�e��
�\36Q��E}�,��_}��@�e�Q���W_K�{��1-����*Q�?3C�A��Y��Q�Ⱦ��(��51�eڜ'���8pH���X%�},7tX,�SzG���)|E��W3ia@XP��mM
Y�"��qLנ��qQ)�����0D�M+k��� �ko��YnN����8\A�@���N�U���+�4��}�����c(�|�cK=\9&橑�ap4F���h��=?|����.QL��@�/��-6��S5��dX�r�-GE���,�ޏ��!��x ��m�wp��V;.�p��?A��FB����L�<`��f��+*<������[���d8�:�豚��I.�v��N�K��V= �����I�G��O	}�I�ⴱ��L��k[�Am��u�-��3`5�!�x�hqmC�	�R=�]S�����d!Q`�"
R�(��"[)w߀vlvL+KJ�ܹt��G~�H��[b�(H���=� ��X*��ǃ`5>��٩�1��I��{o��pC%E`#�!�@8[��狲��Z2N��>׬����fԀ�n�"jyC#��Z�3�bz~|�F�뎓�p�k��P��;%�X!�j2�8�R�x���i�8Ķ�>o�n`T�䗌s�S��4�.gK�B�-^�E�:z�]*�� l-�n�3/Z�jdMG�����U���	��t{�W���AvAe(�|ph�;9��(�rh�'iG�e�Ȣrq5��"��V_���X�F=`��-�-m��Ч��q�3ϣ��8�x�sۉ��^�T��St�Q��M��^Iq[؃�& �����{�B%�=����|���U-s`%���q��"�-O��<�2B�<�YpY-�T���4��P���SlNl���Yh<�g|f6�.��#V��깭��ȕ��S�붐�����x�?ϟy1��أፄ����V3�&Z��&����*�x M�0Bڭs�d�� ��+���`3kƄ��`��[9@w������ϳ�f>�̈�KXlD�*�c�B��d�Wf�,�$X#��.n��J/>iq������#�����:�o����������Q���Pwi�#�P�}̯��~��xC���~R����A�FB����*�R`�c��#���{�w�R�C)�f;�'�JgH�H�+�:`0��$)�Ԃ������ԛ���0��ħ�I-+;2=��˼*p'���s��o�cx%����O�J�(�����Rj	oVNS�?�Ώ �Tv� �X�]|�����	��w���@	�������P�i�*a)����Ձ"UR<��F��.�-�*������7�?	����W�Y=��i����D����
�?J�֗^M��V�L�����H�s?�9c�8���,fq�19���*�œz��v˃�$]��y5�vҎ���-��� �2Ͼ�Pc\�1�����O�7�FY.g>�(�<+$�Ff��2eXPS�&��V}�-������H�퀉_��rsJ���� �方Ne�>�*(��C%4g����& Z?qw�X� I� bo�W�V�(��h�踟e�@R謆��������{�F����v׌�
��m�R(�,Q�gU��I=���a#ޫ��Q���i`��3��#���f� ������!�c�e����d*�.[���w��`⨯�BR;���ɰ�^+�B p�P��Z�i�S4 &�����z�@��s	�uBN��t����<ᰫ�)̆AY��g1���f��D�Q��~ɘ󤨄��;�R�HvG�H����/-TZt/���!r(������}���p��H^���0k�7��D3ڸo�j0�n������ dCEY���O�I�����k�3A6�gb�:6��p@�j�H�Ȣqa��ؐ���.�[��7��ޟ��¨]:�<UdH�%�Itt*)pD�.��Ͽ�3KHs�ʴ��Q��t=��`IcH�O���t=]f��9�g�'�2�P��G$�4�h^�1CB�v�q�Aܜ*�ֿJ-�z6{�4)� ���v!]'͏�U˼��+Xg��gu��*o���#k{�,��u���	�Nn���Rx;)/���{��d��J�}�d��c(��d�dDu��;�� E�T��o�-��iǠ_N�V'Ӻ7�!7�������QoM 3��)�Kp�d��I~�mb|�Ƀҷ��j�s��Y~��3:=	ƨ�%��~�٩-�V��hdᔆ����w�1�ro+��6���	B�ʛ���W�Om�����ey����*�{�;�ޜY $J�j��X�Ñ���E���	�y�_n�[�<�z/W�b�ӈ��$zn�X��6���۝g��메��5�}M^W5���(6ȁ��PI�B��d��F��;������.pn��xu�!��� �Y���7�M�R`=��wڙ��>��:�����^��i?o��S@�Fi�?�{�ʏ�7W	�m�ma��*����R���bHWV�1A�-�硵I���)��d�z̴V����8�Ie6�<}&I���Chr} ��4V�7�@l"
�[��<#���Z38�K.*�wG~`���B;��&��}M�b�� ��U7S��hl�~b����7L3Y]�-z� b�1O,��n0�a]��dVҹ���̳��� \�w��x7���ZN��d�a�3%�'�;�Y=��,,�,�#�-����K\|��R�����=��������S�Y�yP��L~֬�����:�����4����W�����e�N%�P@��E����_Ys�e��5X����k'i�ݖZ��X��%�	���=�_�q!z椼Ș������y�y^�C70�הG����B!2c^�m�&��̊����^�s^��+ɫ[�Nc�M:4�� (�U۹���E.qot]��VM$��F�3t�5��6R�w�p�<~�T���F�XC���ޝ n5��|�Y��ᚹ[�3��'W�]X�T$����@��-⡓^��>W]��ɻ{�G��P���p#�Ԥ�����ɨ6�pl���ٕ{���P�W�d���kj��ll����ϊ릥�ƅ�����L|�-,�]sW<�c�>_~��?b�t���8�L��!�|
vɁ�7!W.�b�����Q:2ø���1+��^*�<��o5�ӷ�8�d��2&��)oo���̧)sS���lS���^��hq���o�Q���-��뗶;���A�}4��Ųސ6��5���� �>�Nk�lz�~L�=eR�����?آ�6�!)d�>������fPt\�x.é��~����dt����%�;R�F��X���'@X#f����Ɖ6%���+���ol��PV�|{z�
 ���D9z�f宕�8��	yDC������gn=�ge��P��S.��݉RBƉ3��2F�B���+\L6�^n���f
��T��B%�kg��]���3r=�Ò{��nhRn�o �L5�3�A0<�h��<C��a��<���<DUm�����~����CͶ��ρ�~']�P���+3��z��P��Rˬ�^DI�'��e�R�+0ΣlG��O*��YH��Ɇ��Qk��jj"��oZ����?��l�$�u`}��\v�q�U��ܓ�z���{��>��(%Jx�z��0I:kd�)>��c�<��>Wn� 9�%0� � I�0'��];`9���E��:��~�	��X�6�m�kM��7� �^��6�5!"o�b�5X�~�N�ɢ�Fc�MS豾�K�����Q����Д�Uz�OjW��d2|z%��)#�
�
�Ϭ�̓�����j7�����P+�����γ�I#�>}(�s,:�Ո��Vr�Amϐb��|�����LU0��MI���7fq���N#5p�"��:߮����	1�����ё��������Ux�qW/���}K)x�4D]�"v�|}�}�p�E����-bg����$���[������.�؆�jJ�]�͘��v7��g�-�ب~;��e
������A9��֣�HS�[{g{��xۄ^;�����[\3� U � `W_n(�b����G�qT���R��8^���? a�d��_�!�O7���5m��H���=��}��:��ϲ& �0��J��	��Z�Z\|���5�a�g �/3ấծQy��.;֯
���1���-���__dS�}�����SBS�k?2՘[�Y�/��õQ��i��U��Z�[��M�ŧ��t�{21^NT�L�h�үO�'�'=�/�@�]�	�	��':��|�T�d��f-v��?�m�Z�8ٌ����B�mtf���-���%q�
���7�(�[m�4mD��vCu.�K�����)�Q�E`O�+���
3ԇ�M]�4�ꙫL�[�\�B��3����t�C�U33��Pq��y�����=f��P���[�R�H!���gR�-��P��ry�b��Ѯ���4�E�]�{з�RRh��3
�;�����	��2���{�K�KN:�\��4�0%�[�A�~-X��W3� �Hb$�����d-�	����9�~��R��6�\j��[>t�v�ϩ5%�e#����;}�T�����fH���lFNbR���޵�o��3��?@/3VY9]��E1�,��ڞ�VmB�/�^�*�(��iZ���p�~X߳��e~��i��p��ї�(!hA��ע�g�"�羊sT��Q��*�Š/�t�<'��;��d����V�1J��g�a	����S��"�j�Q�������ɘrrP<\y7��/?�k�e�����D�FR�U���\EO�_i���B���nBEy�6OE˰խ�=����P�m3��ԧ����k���?��Wj����ˠi��D�-�M^Q{�i��J
g
5�F�bc~䳃�f�D:�o�:,�`j�=�)H:A�z���
�߅	��V��_��	��q�l��Ǧda�_+Ҋ˴��)�Nx)]���ƕ�t�h��hb	_~^�~rto�@T1=�u:vӮ:�R~���:-�	T�sߟ�����L,�_hl����\6�#��^�(|Z'7��^:��������Ǹ\6��T$���w��KV�9���6a�jL���t�n������Ƀ@�,���v�sO�;z����دn6=�z�(-�?��.���^�t��NuW5��W�Pِ����������{��Cˉ !	2�k��1c �"r���R1	���а����8�������HS�"֫�7�޷S+.3L�e�alfn.����G�g+��d�Pn'�&|������Dߖ��"��C�=9\
���AV������3K+�	�0����I�w�U�\t8v�I'����+�h�U�����>�5N�̈́I�Ɠ�� C��xn�QYa��m<��<���Q��*f�Me9
'X/P�ɹ(A�R��#�E(����u�i{�V�#��u�D�Y�W��ʞC�I���R*N*}�4;��w�ٰq�0^�{�o9���W��j��J���B��R��n��(���G&1��.����F���3�^�'�"O���{��&��ӛv?w�DO��;�Ǝ��5ý��|-��+:'�0_�f��N�Ȯ���!c  �o� |������S�\6���Ul^��v���!�*�D�`��(s��A��q�?�ɥ ��C��;��O�_V�jbb`y�\���� �Ƙ��Q�R�hhSj�#f����/&T������f��@N�l2���zk��@eCE�{�ZT#^�"���P�"~��q��.|:��T��X�`d�N�7u��*����p�Uyʽ�³���B�0嵙p��Q+���2�׍�zA�:��%q|����Qiv�I��k5,bM��15COA�󡜲�0x��q,���4
>��Jf�Z0.��a��Y�B�y.{#��^?����~����ϒ� _	�r�%�j�������!s��x^,�}
^<vZ�k
@�@+[��zip��$�4=#��Wp�X?	R�X�䛀a���;鬬�H����k)��'լDS�
BYA}�K� �ƚc���uI7wmZ���[��_���ծ�p^��/�k���Y�(`Ts5��űeh�a�|6߿�J����E�C^����I+JI�O�bl�rn�iT��˥w�!��q� m<� �4�{�`o��ݒ�����韟���Z�2rci��f�g��EkX|���ղ�ֿ�i��$�G�'T�p�]�X1���R���o�
��x�%5����Z���॥|<�U;-�G��~-[L��D�gެ+�"�A�VJ���T�aoЪ�LL3�^����������=���h�������fR��p \,�<g��zj��/�Z~�)[k��#o��{9�s��k��|���J�+띲�ec���
kO�QB|bc�w��
�{����xQ+����}���6��U���k�[жNZ��kBZ4�7���̈́}���X�E�c�_t[0j�(�@\X��x�[�*$�z�R#����&s>l�fg~�]��a��x�Q�! ��o��ɝG�αO~u�a�Qb�LY��&����K��Ъt��0x�.�N��0ȇ�;n�o����51b�p�at:�qG��{�K1"���ϗ8��?���MqI2�J�+G]�Б��F��R�~6*���9��:&;.�0��o۟�ː)7��:�ߨTFە��>>�K��+S��'��Kx�E�K����T�ʒ���N7�&p@2�^q�ؒM����٤�D�A�ߛ�Àʺ� �r�a�{;֧��=VS�wl����b�AM��h��*+p� �3 �����+ؕ�%�_�al� fr6����q�T%p?	 ���5sb^i���@��q���m��z
�0�AJ����ƽ��_�%Jm�{�٧=�"א��D�|0Q"��W4���K�bHU��o��/c�JGJ��bW����S</M��^�jt���)�a�z �fd'�t��j����,ܯWXHs��D�F�;�u��}�k�]�Zm7`���)����;9{xHz[���bs�����:��+��I8p<�s]j�Ý�������q�L�a*�P�Hl�iَ��A�W��*���'9�@��K?M�q��붗<?q�7��220T�0��w<W�=��-��l���),��ʒ�[��=5�4�F��e�^��h��8�����	9Z�&2�LmE��e����B�y�ɝ.���ЃȀv�g�c�>^+��1D�px���b�	x\)v��e��u����r|��߈�2�?��\��z�T-[[;�!^�����$#���h�v"��<Le��iO��S���l�w��;�}���^xX�� o�$IQ@2�V���W*,3���[��w2 ݇��j�	�2[�;�� /��)"���z��[�i o�8���߲��3.�#rr�@A}�l�ap��T�T4mY��aJ���ʹ�?Я�����C;�:N����	6O�)� }�ާFI�:{>��|�����DMsL�*���?.�h����_���b|1���2���R�6�6E>�� ��H���Mў�;�.c��N
�(�T��Qf*�&ZZL��7&�E��;r�G����^B�.�"���v�;#�<EAC��Ȧ�JKҴ��]2��#�Qw§r�Á|IS���}Mx�W+��u��*�Vn����N�� w���C��hx��/8�X]xz�F��N�H�Wz����		}`���Ȣ��N[Wt�.���n�k>a�M��J��_�R�벞���[O2C�E�{�d������0���a���G�Æ��4
�4����8�jno�d�tUez$Ih>����Jʢa�� /х�╌�w6�����h�3�hNH�gҤe�杭g�]�\��϶�u�c!�s���m=�Pli�g㆐l!���AE��W'A%���~8����`��9�$��o�^�6^���ώ�O�A-<���R��_D}���>��(I�vFWL�PC�U�	�a�����`4іU���� q���K֭�|����Hi<��r�T�dI$c��;�mw.�����s��tK�1[����e7d�`�u#�$��Ñ��d�}���q �ڟ_�8�.�\�Ї����/;ЪhZ�R1נ��|-S��ձ�0���2����=&�<���
�G����9V�l/_rE��g�23��r��j��	m�'�$Y�\Q_�Xq_�"'<��ư�B7�f�4t�pV��rJ>��;��A��'	}#B��>�ާ�d~��o�Y��v�A��躟��7���9\�`�:�jH2���%�<pa(q2W�'p ���u�!l��UxC5d ��'��@5��,�h���LU��;��V,U� �9 T�B��^�8_kWH�G�e�\U�G�s�&t��.�I���n��\����#Tސ�y�?��OA�Cw9^���H��W��lȹ{x���O	�]j��Ռ�֕��+o�y��V��t(��,@��ښ�1iW�艛��ĒT�Q�@D�ǒ#`���6>���h ���G��ef���^.j�ǫ�G'D�Sb����V���*�Cw�"x�$��/��a��Q�sѰ�[:���+�vG�'v� &��X��bm۞;�M����
6
�')iٶ�m�k� �eP�̯a�n��Y����5�Q�L�R�XXǈX��w2�"��L�A�<�̀&��?*��t��3�>��p_�n����
�S�X|��eM��O�S[Xx��s��g�Y�IA��p�b7���s6��Rf*��B.�\��w��}2�`6�F �
� <<~XIu�V��������HV+�l �?�q1\�!R�7D�	O�c�f�h|\h� �>������܊8����i����j�+��G#��W�:��_
J_W����!��3�v�G5�H��l�Ǩ�$
E�4~ޓ�%�^��n�.0h���+�'�+5-`����6"M�0����ӎw��L�����"B�ƺ_@8��1]�?c}�J�<�̭*�̠�����gFq/u�1��'��]�kHS��Uo���R�l3>ѱ�"��8[�������n7���i����Ne��Ў�c��X8���3%�ǻvF�&w��{DV��~rQNB����6���]c¹�b�B��'/�ٵ?�$�\.0f�KYP��wΈ�^�|�J�q#�L�,)�~�"�#��ff*?��O܄���z�����0
��d%�c��]�[3��s���4��o�-¸3�`��$�aVF�B'�;6�}�f�KS~��7U�d�&X�K����Ѥ�6�l�d��r�ڏ@�&�&W��z���
? �5I���S UΧXŕ��3����+�?�IK�tb��?4ƿJ��~ѐ�8�?M�/@:�����nnm�4�HP���A�P���zhOl��Ò�e#��>O�{5_Spt`џ�
�æ[oJb�F�<Xۆq�{�`J�}cj{��]C�Z\p����-��ɠ������ٔD\��Ƶ$�1�u��+�з<�^�ȶhXeg��C������[$=+��	��?�Z@���ҵ�^^XJ�"�FB��56�bB~|������]As��h��Oxf	l%��7��&q!�_&�E3#�V�n#=i�eM3��(�U�z~$�S�΄�(@�ms�3T��k'�;�M_SԾ�����1昖r�L!t�|*�u�L�)����WQ�
&��A�!^e(����v�{Z��k�P��ER��[��l�g?G*]��z���>��yT9��zkY��u�	BDW��_yML8Ʊ��=,��e��-�<�����pO����Ee4Cx¾K�
�ύf����O5�O�B3Q�A�o�Kw�AsB��?�j�7�w��2�
�DJ�57���:� ]�i�� �w����/߮����kwx��M�n|MԸ3� �M�᭚���Y�O�R���l��f�5_'
�e���zԚ"2���N�u7��[N��D��^ٸ��,����˭��l��#�ez=����j���S6_��\Wڞ� (������&�,��-zĢZ�z�R���X��dx8~+36�T���w� 
�
�뫧��:���uwN�i��+�hȳob{��0�<��P���\��WjA��g���ⰇG��
(�n
.�M�}y[=-���L�
x�1���*���
�ݏ���] ��=fĢ�q���0h�)���e�[�.Y�LK��bV4������X[�?���φ.�n[-����[���Q�xg ����PHڇ�'|kKvv�@=�3v6�x��Y�jF�3�xN�D��3^5��P�W�U��?�����߆a�ܻ��B���×�^��NN�Z!��>N6l@lt��y���{41 }N�X��w�?�G��'	.�7�;N��޻���9�:��]%��l2+�A�⵮ :\� y��������1c�;�$�=���
���������5:R�WL��N�9 �%Eo���ԻL����t�����m�tZQ�����®� x�q���3��_ј�]5�����p�������6���Ƭ}�����L$�!�����J��8��h��X޶�za:ߤ���g��!�����t����{a��6c�����(Iͻ�w�_z���"9+0��Qh�+������i��6bܽ_n�E��qpzI��m���僋�%ƴt#�-Y*�\���^�&��²g:hC�}_�I�A�jn"K��"'�C7s�b ��vw$@��)f�ݙ���i���\�]�t��Ҿ������n�}����<���#o�|'zY��rY�˱�TAR�2��D�g��9O�%q�-��F�$�U8��0PTH���=���<��c���[ɉqH��w	�膪Y`�^���²��X�Z���/��q�Zj��&�6�����.��6:�!-��y4;b�t%X�ȁ:?�d }�N�7�D��O	�]%X����џ&)2�:��LC�V������s].t}��^r|�"�؛5�楝w+"V�$��ut��j��G���ހ���qfF��vޢ�#�j�	Y��@���A�5�A�o��+�H~�2�����q�)�.�V5�)�Z�6H��n��?6�S��_�`�L���$�����=�B��K;����B뷞��(y$D���ԧ�О?�>���`�"�'����e^Z��:%�~P��ehu1�!{5@:�'��������
�"��V���	��a�ɸ���[�gO���<����,�	 g���g�[o��565˝��6�{	�~ߺ��;��(nBK�������7q<�rH��3���M~9^���.�n�n�E�Mk�I��:7���=x�y���q� �/�i���(��*��eE��b��䌰�L���!��h�>�Q�D���1���%q��
�^�ʤ�.�5�SC�eE<���̴k�H�h�XNK�߾ֺ_��Z�6��~�"u��"��zJ{��q�oh6)�-#G��f���b8~��
�^�j�&v�*` ���/�[�v�����H*9��r�H�~W�E�8~bF�9-zl�cG�⠕�ѫ���Qș��A�m|��^�<���m`;�1W�oAd��̓�<s��6:kX������=m�I9����͌�Z�`��3���-�=K]cLo%Uǐ���^l�����X�tc/�Țа����Y���"�u�:-e�x`�*�X�q��k���-6�X�D��2�`:�"!��%�����)>`�w�o	���alI���%�2�Gl78����$���]��`�o_�ō��v�Õz�G%�J�(VBC9)�mX88,#rp[ ��5\j�7��*���u�w�.��m��`}~\�B�h��4�.ej�ʱ���;�VD�f;��)�"���;��24ή>.9|� S��^VQn�qd�[�sE��E�z8v��2��	���i�i�<������b��bf��Ȥ_���I�L��
�	�M��� ���A1%BY�X`?d��c���`FԾ�!��ʵ=��������1��Kl�T�9Y�LV5���O=Cњ�֝�'zY�>E��5��F4�n�hϷd_�|���N�=s0�(�n�}��y~ó0�{-nS�&;�ت+����� 3�FYY�'J�y�jE�<�t�ˬ6ԄW�/�2���m��a�����_����5�a�p"��]�f�+0�S��JP��ע�O�l2�L�9ɺ:��/�*#�Xɝi�m+�R��S�b�.&��i �*!����b�p���k� e�U}��"��?c� 4�2}֩���5hq)�lE��������E �+7�>���|6S�;	M*����c���D���w�0��0����˝�cݻ����՝[��=W^v�����	ڛ�}$����$����n��`�gӺ@X��Gn��T.,Dx� ��$:�Ӆ��*1��xa��D�Y1Ar��b �3��]P���;X��*k)R�4����O���x�4����Tt���D��q�R���]NA�P��
]�-�s�.�iI���3�?5eP�i�5�՘��b�bW��`�����zbC��x�W���6l��[�'B.M�bgխ�0�0F�p��}����7O��=>��x����UĘ���QKo]�M��h'����`�M���) 7�X�p�{��j-�?�d�������e��(�4��ד�^Up�p'���Q��0�����4C�1�n��=mN�n#C	����}��w>�j�) 8�t�U�E�#�Qм���p���
7���]і냤;��a�������+��Хލ�l0h���3[���Coڑ=�R�70�yi%|��51��P�~8�jp���7��=�uH�:g���Ɏl@���x6���\���JpJ݅ �]���i4�E���x����=+��)��2�t��m/i���f ��N��
��II���s&Gg��Ò���ORf����I[��W�5�C��β�g $h�a���C:Fv���Xq����~�������zQ"��s����sD�"�l���V��6���C����h���>n���ײ�9"�C�`ZO��!�Y<����<w���9{�q�K�����>+[A	���L �+�`�1p�#�7-U��(36{�d��)ڴ��!�I��Y�wk�7ԏ6������ȝ����D�k7�?�F��pu��/R��j��$Şc9��I��btaY��k�u:F3�Y�vm����c:�q\f�ŏ�9��I7��*�$�h��<�}<j�-����r�a^���ї{����� �KKh|��1�'���[44��ǎ�*��F6}���M��X�>��X�?Y���t�[.]��Dch������S2�;4���_8"��9j9?T�jE��*7�l�͘�0J��ü}d�D�V9������'�x˟�2
Z(Α��OD�q�^��@��A�5X�v�_+ɖ��6A͘~ӑ���PNq0�FbG�]�f"��5{	��Z|�Do�Ci�!����cl��9&?#ϒy����:�`���A LaԎb��ݐ�u�9�_:A���"o�o����&.3��_���q�W�sj�?�����`���wW��eƚ1v\H�Wp��dsB���4~�q� �$?��X�խo钨��-��C�HU�?������'Wo�;Y�T'�23}L)�y�~Hk��tk���o��\X��$�Ϻ~!��I֚.�O��_Ȣe����_��g��M��3�n�GtN_����@�od�h�7��7��|~R�=�"��W���l�%4��v&���v.tunV����4X�8�=η�c�a�]1�x�sc�����Ұ�`�A&�;rG/��'�ۭ�]+Ae����G��l�-ǌ�}*g���tDT+�֫Ig0k;]]�W�ܖ���^%�$t�tzk(əe��5j��	Ͱ�5�N��#�UQ&Jj�d����ӃH~ʃwh�p1�Lnw@Ɍ`4Y���+�pm�~���x���a���>D�&��j��G>�i�O�~�v�S��pcY�F��nͫ�b񙡌�W�!-V�J���I? ���>%�]�� [[���nA& �xS��А�H��*��]�ȞBȃl��	���
���'v��˅> ���t���T��w#����׫@�ˑ�d�B�;��!�-�b9j�����"B�=j�� @����lݔ��%��1d�.Kێ��f|�j��td8L� ��� ���J��}���2.�b~��N%�i-�x#G�H{���F�H��pZ G���0<4�Mz�/����#�C���LȎ,�`���l��Mx8M�B�n�z�g�j �["��Oo}���aH�
U�DJ��τ;�����WB�K��]�mp}���`�X!�Q��]#=��M�=���:R�}?�D�rm/�t�v%BQ���|G���3��ஐ8OjaP�">�.�s���g!�X� �����,G�M6~�'�TD��M���PlM@����nS��C#z��e�w �+.\�c|�P{��^��.%�ME�a�ݤQ�
�B�.�g�s� K�ǞR�k	L;��7Z2�r!N��4�ZMv�ug���0䈆<e8�A.�������v���N��~��q��__����	~�%�0��A���dA�`ǲk��]�T6E8Օ�q�n��"sMH�[5�F��1�w��!�%�k[�.S_�x3�?�zp��8��N�B�j=�__S�Y�ϙ�7��NA}�l�X֒ 
.������uc���5�Ef_��`ر$U8�ޚq\D�M�9�����8ȹ��8�)�]��h̚����a��Jg��c����	s&�ţ�%��s����%+	�� �Ӆ9�튟Ð��1æNI
�=��Y=��`�M/�e�vuw�[e�5��[g��&�.;���M��h��x+Y����C�DS&����B�����T[� ���	����%�oi��E����En���V�ڥ~�WY<"�G�{Ә`���B6�k��Z�
]YWZQ����(H5�į�,�"5m?+<��j��o��%A������S~!�Ϝ=�²���hǮ6)�# K�ޔ�4<!X�}RM�L\jG�$�T���\�����-�o���vg7>q>�^8Na����0��6NqOnriD��# �ˉ���qkc���.Ĩ��(��� 9As�����
 g����>'�rJ�7$RE#�:�OiA��i�o�s1$���7t��d�{�`1 s��`֟�&��ru�}{oB�RӀj�VSxXOm��|A��<���ΐ2zz�Z�m������Gy�lp&']�	
��;���[����+5�87�t�2C���,����:��9ʕ�c���Ǵ�}h�zP0��{ǬiQ��H�}�m�y=�Ԝ�̣�3�T��kK�ժZ%+o����r�v�0�볚�wծq��@��vzz���<���H�	QT6cd9�41}�D)����+�"�:z�ڳ.�	�S�-h��˃.2$���X5��&���9brg"[��%&h������#�א��^)�_=|S��?ư��1Z��]�o{�T� ݐ�u��;rv�b8N�
\�M��`���L���)?�y;'y�zٗbd��ɣߘ�r�y+5��޸�����T�� ��*F3�N�|ar�d��cʆ���۲�:�EA��K9c�K�p+���d�/65*��08�w��	H�e�f���P�)�@�l^��ś﨟fyzkS�~�	�;},��q�EΆD]�k� E,x�:'-�,�����8���:1��^L[��՗�y?�H����8y�aꞷ'�ӽ��wy�)rE��rh�YG-��-홊}�\���������f�۟f�y����r��p1�)���=%EdA���'����'���t�N�Ȋ
�٨)Bl�rݱt�����7In�r=U3�K~�9X� �;���I �f��'w�R ?��s�	砺�LS��d|�D�%K�����8x� ༫�%����Re9ن
�a\MO����y�e�r���|��10O�.F����ֻ)MtCm���`si�ox���{_̯��;���3��늆?Z�B�@Z	xѡI�m
�rܺ4�$��B|l*���ۚN
w����:�5V��M72iӞ�?�dX����|8o�&�a��AaɓO�];%u�v�6�����K�8����t}!�5��\���ݤ�`CL�Z�.����I��tU?ԛ)FJ�ܲj�2Ol�n��źcb� �=SL'�~/K��0?�=�oz "�A@:���_�U���i�ȕK��T@�� qH1轓���l#>Z�/����@�32F%�]/\�X�:���}�3$o�}4�U�g,�v��%�Bd�/���,��Ss����v��fp�h1�M�Cꥰĥ�Pw�`��9���+��� ����iY��0g���a�bSbČ�w��fƿ���J�&>��Qu��]52��u���rC�v�EEO�cD��(�>�_q�s��Ǒ�j=�8�><ФQ�5'�^����SM�;k�=(��nWk�eV4�ˇ�h���7���J�כOA��h�t��C�D��72�.ѽ֟g���-����rѹ1�K�h�@���Uǲ��M �x ����`#����t�ӎ5ܗn�Y��̢+�~H�,�O}���
,\i��Ϊ�0K�6	�"�Y�E�;��mEj��+��l��^��G����� 3� ��U���#	;(
�{����Ȼr��ؕ�{(I
�o)���$D�1�kz�KKrD�b��@��B�����76H]\0�RibJ�ɨ���csG�v�W�zOU0j̮� :��xE�s��&����������ﱞp�E���WЅ��1��L!ꚫ.Q���+a��LyjY�묓�N���Ra�("8n�vqſ���K��w	��i͋&�sA���]��2iҳ\
�I���}�	���85��Ǹ�̒y�I����\� �F��!�M�0��[��J=b�*O���1��Z�IH�\{&/S^t#�@cu��`b�̥^��9��VY�eu������g%3K�±�e�I�.�u�}���OS@�/3?r�r��
����l�	ī�4��}��-�\'c��T����b|K��>��T�ddP�F-Y�\����y���1������L��@Bp8�i|�V$Yc�Wqk�	���(htIIQU�P�ƹ���K�u��g�����"	&8ʶ,� �k7�k��z`��l3ǟ�OS��t�	.�I�����&���W�q�)���P�j�k�\��-讼sW�=C����+�1��8V��o4h �R�����oGe�JL����N����Lr]a� w#:i�=��&[���5�=�{�VO]���e���:�	�juC@�Q����q�LdT�.�2&��`�钒��Jᢊ_J�x�=D����f40�]!*�H�o�u��5:�4P�)�ӳ�flY]���O���#�ZԞZM�b~~��{47�/��I��ßeɄN�;}4�%&.fd MZ�Y�%2G1қ"D�i4up�A�k�&	K҄Ҝ~�F[7�~�NY�ML+.�4��;o=S�p�SɅ��)�~��^���d|8J}@��p.F��fkoVg&���W�-�D��Lǽ�Ե�~ XO��,�'�������ey��P `\O]}��:\���\( Z�͹ zd����T��$b"���LY�3�b,Z]`�|�ߊ��h(�,�6�ȓ��L<��I�������2v���6 �Y��GP���nRB���>�,wm �_=h���E�oӗ"��Ob�s"�Y�D&'��N���8�PZZ�*�B�{��JE�����`�݀ȗk�'U���
"�F��_(t��r��2��8D�J���i(�:`x+��2B��G7� �J�t����:Hf�8�3�&�|E_^S�D�^��s2����o�8���j��e�u[�/2�uM[�L�sDے��z�WF���=�!4��߰8��F���-Y�����kk�m?s�`?к��
?oZGU�-T֒-�k�x�S�pCQ��[��s���T�#M�:�4�Kf�YN��t9s���2JȊ�������).��#�A;f�S,?n��ДL�H�H�l�p,��B	�M�
[�^�hV�-���t�\m� ���+7�1�N
�.�KO[VPƣ)���x�77��:�D���ʖͱ�~pn�󻅇2q�E1碹��"���0����%VS�L$F�E�b�=�AxQAw{]���H���tV^*��L&=.�@i��@�ɯ]��R��^L)�r�8(6kG����N���`�Ok����~�da� ���y/xH5Y[Dv�x��湟�A�.�JV���k-u��֤a^���H ���X�5�¼-�uL��.8t=���Vv��V��L�>�t���R�Z��椄1�H��.&%�I�MHU �����ý��u�U��k�c:N�!9_�G������3�T���gG�� p�oF#x�t� �ͫ�*�t�� ��+bO�dN:3�5dS'2�g�5���Jx3:$x��A��>Sє��F+}�pw��L{�6�S��[�9HR.�hό��(i��@�Ң�������mY"g���r�,���،Z9�)婩5��(�ʰ�.*�ЩBF�0�:E�f�h]L�l�c�I����7�}2 {�EY�١�o�#W:��B$]q��<���E}�	B�U�L�5A̫�w� �W������JGv߹����Y�=d\#Ԯ���Le�=f���!xB�y�tg/�
;��R�JEd�H�aa����Q?� r�Z�yg m�������f='��
��rl̔3hЈI����q(�!B���/�c�Y���B�C����5��s�CB,� d�mc��U'�G���ҁ����:��V�a!n�8�������}s���g-3奔o�?�,���=\��L�ѯl]��>�}���Xgc�"f�%m����-}�/\�:7���M�C��=��U'��抉U�����
���my7~�8}�Ҍ߻*a���1����Y/�d�OR1(�h3=u��]��jT��$�c���}vMbޕ��j��X���[g7�ɲz0�A���d�cJ�,�+/�a�{�܀�=^Y��O?�2����1N��J��e��_.;��O���y������C��������G�bm���0o���K��`/����uC�H�H�+�,0�� ~68^��%wV�����!�=�����T��_el1b2������~/� �c�Ĕ�y�'8������Oړ����B��z�'@l߲�����)K�
qF��J���Og���Rǔ�ǌ�nDWE*�ѓ]��X���u�	���g����ﲢ���[�;y�׈Wt?X�E�Y�.��C�q+yNd=^X���sO�M*X�.��vh�թ1V�� ��h64���������5laJ���eMo�����6򀷂��uժJ��1�&��_�"Щ���-_?1:�'�4ȇ�=�b�>>��}�E�Gq�=��y���R=��A�z��T�[z�J��
5Y30<�:�	-C��D51n;���6}A�t�<�tml*F�r>@��a]��%�[[��j�6��@k�+[�сvܱ��T�b����~�N�yN9#�
/|�P>�I\FlM�!#�l.���W�G�X����@Wo�N���Z�������_k�V#���E�J��Z
m���o�IGr�O0zx(�T͉D?f�y���J�7�D��K�/{�o���Q���e��&ϖ���&C�6`R�OZ��(zS5|���1��NP���%-��KO�$M2e�*4ћ�<9��,���wx�(�>�^bS�wv��͚G3��R%,�tw��.,�cB���t�P�m�g���e�-�v�N� 
���O9lS�/v<�{0>yS��`��=21���
��p���@�9{��$��2�4|[���B�9�p������V3�Ŏ��$�hƅ�������IU�V{�Je�Tѭ �~d,�Q���<�dDr3G~$�܍�5�!���G7#:��l��ĺ��|>Yɗ�N=ɀx����ӗn�Ձ��o�	�V���}T+,�|w� ]��a��,�IGkm7�Xplš�O�U;�,�N��4��g����rId^%P�h�6h�T3<ja�Ɔzf衎�8�>\J��J�����H�i�E��|U�G$��9��_1sXM��A�ܮ�9�h��@k��桷s>������O�L��@l����/��gU���VD"��,\�޷ʲys�xK]����Öf�C	���r� f3�r�K�t��c��)p{rJ��|��q�Y-q-|�De7��m�3����M�9~QiIﲲ7?U]ϮſK��z/$Ӻ�h��@�h6�UOo�bx�|_8K�ڠ61��N� A]�thy��m͆�����0er3���5jN�=�_����|^�S*K�[ez鑌� ��L�򇾲�c�rԺ�l���"�a�Е�S(��Q���7�S��S�q�ٝ��]��gkz�P%�����ٽwo<F�lٵ*2�F����CL���ĵN�`�[q�ߖU�4��k�_���w�4��HȇL�$aN<�XR
'�.|�y爠���U�.c6���o�x@t�K�to�Q��J:($�z�s��� � :�r��&ח�ӎ,wa � ��bD��a]gg��ߪh_/�Lq�0O�L���:�we��rs�`o�fU�m�(dF�+"�XHޕl#�)Е�FbJ��A�q⇦��W��$�G�]��H*�ɚ�;�p��l0��(AM2a��+��ua�fI�{�B�]En㜑Z��gƎ"�>'���
������b�� n��M?��� �hu��	:��7��)G�F7�������+^̫���̲�������d����F�]U<�$���_�(,�q?ʮ�^��
T�N�,uU�+V��A�M�6�Rf�c��!㐖��M��}L��6n�������GT��~$"��ږ��0UF?9���O߾1�Aw="�M{/���t�T�"sd(V�r�	c (�z'���\�9�6���8X�;��r�-�Z���� n<�e.�b�R�B�f0t~�N`Œ��+�!���|�$赜8�y�M�T�(B�'�k�4PA�M��Y�<'��h$�T70e�H��ne��ʧ�20"& �v��fa��r��T/q ?�խ>����m�j!�� ���{Ty,��ͮ#��=��+?k�[cZ{4��p6�>��ް_�BGz���d�aYט;�ٿ5����PT|T����`ϲ��q���2R]��q����Q�.��*��fo�Z�}��V0sN�4�B�)�4v��0�r^��8ⓞ(4���H���އþU�'dck0�c(v?M�6�rw4�w�"���	�V�u��*�]��6#R�[�`ƯBF�������f5JؿH|�r�7/�,}dtAJ��dA8wx�`8�ɫ3�w�ʵ���ۆ��*4��E�C�Ϊ��Fi�.��('��vs�{�+������k�6��A��U�!�,����(]/Y�y���ḉE��Ĉ��rg$�WQ��dhp���u	��s7�0�w���^�d�Qt�W6:���F�ýz���m�͆�����!���f��3�}Y��>�?�h��`d!O{[h�n}���:RƉ�����-l&��m�?���[:A~J�����2�����B�[����Y��%�ћQ�9?�ʘ�����&T��p4��P-0�7��<1h��L�nP娛 �2�O����n�>I�$pX��x�ƙ�m(�E��l��9��F�]�dݽ8��g�
-��5�ǂs1o_Ρ&k�p��ǰ:	�=� �=a��cHg��U�ӳ&�Q��Nl)0��*sw���՛�}KR�u~�U�j��y�qyw�]�ѐe����<��>u���Rq�E�ĝ6H1h
�"ׅ�D�=�#(�����"�и�fDTA��'��'��{�p�R8sˉ�����M��=�
�~P��5+����ȱZa� +�'������K���
M��q9�Xu,gi�J��Al-c�5�r���z�G	�nXS��u}b�$��c��Tr�[�<k���/�zB) ��&}r�Y���b���C�6�Z�iG��_�5�;w�	1�P���7(»��z1�H:��b�O4�?M=Wa�!��X�C�M��D�g��3i8��we[]��-_S��g7��(����t����n��쨛���Ip��Q�UZ�����|��6�l%�;5{��琐�d�֟�4[di6P���������ch�f&��Ms��4���I�:1�0��l'�}����9��c�>�k�/�[����&1龓��9]7p�{�E��pK+ퟖ�^0G��Z��.t{�[.^N�=���hK��HC�RG�|����r�:�׷�]�v��ژ�.�J�^��˪O���ϐ��LU�����e�e�����q|hT�i�C&s� �yN���+���5/�*xF���ۃ�6O����HT���6Xbr�Q�:�O���mg�ۿ�<EmM��lՉox�<�Kk��ՒD��h�HNFP�<���%!5Jo����;�jlL���pg�2���G��+�-o����[�٫ݠ���$|����)��Z��]�4ך�:�cuP��-�Z�P���b�;r'�/I�����,�I�)u�Jߨ�ڈ�d�3�
3�����r��G=����q%d[�,(a�Ub����ܿM�4#�	h���U�_Oi���j�E<gj`�x,�A�	�%0X\�9�
-�e�捪�pN��c��n��*VW��m�\�k��2��@+�p�"bl��u��
)����Z+��l�A�qǄ�^��KP�{k��	+�K�3���N���wv���K����ܨW�����
w��U�bɤ�n��/�?�0���
z���7�� ��:B���9ƣ���e��B��"~�9?K7��W�|B���۶wK�0lA�?@+���a|Ѣy��n�twtr��j�1�5��ŔN���\�s�� ��jn�jG Ǜ�������K|�	�ˈ�|��Y2����FD(|. ��Z�6������"H�a���*������^�cPo��������	�ې�S��J�ޙP��\f����M��^�VX4�
��_�D,(�0y�����G�u^�X\�B'!)?��{&�Q����b�q�c��$�&ԝ�Qf��{�;�]Q��|������O�'��}8F��9>b���� 0�yi��*o��.��=ɿ���#�� ��fex-�
h�v�p$>1:Ҹ�c�f�G0���B������զ�ıFa-��ǯ����N��@�+Ő�0'*�vɒ����^�*(�J����ת%���t�wzjή%��;��YD��I} ɋR�4�/�0��Uy+�i����܌�/*�jd��Ɣ��Y�'�B�_11[��L<Y������b���#�n�Ҫ�O����S�];Ӧh���2r�s��j���ͪ)�TуǾ=��]�@?��鯩��i��D<�4���6��^~U�`ͯ
����M�G(��*Y�t&"�
�n �s�B�,�s(w�ae��N �TЅc��.���q8(Ƌ`��*���x�ф�T�D;uݮv|�"���\��k+c��� �)G�s8��J���j�A)�����,�5Kv2Mc$J\Gxt�3iJ)O��9��¨��#Ò�軳A����}7���e�O��F��{���Z����w޷�6��^>!F�F����O�A6p�'/�L�z�Lm���Sբ��U��zt �H�4r		.>ϳ���s���C�h����r��d[�u�����.ܧ)�ڗ]�z��t��/�Fb9h@S&��e]g:W�3�W��T��8-�[��kx��}Ri�Ȉ�O
7@��m,�{�25���L�H]��S�_V	U �Դ@�������`Ω�V23Y�ǽw���Y���N.�/DFp����v�<�O���Y�_�x���`�o����Y*�����'�{z͹�f�/~>�~�ZKQHjO2���w�	�c�irl���!����_vH����ŁQ��s(ȹ����?���^�i	=��9Ll  ���YI\�4�R'�U��G������YG֓��L�y�Gj\A�:��������[��{m�� ���EĤ�}�8�����D[b�tZ��wW�I��[��W�_�K�/:
M<Ň{�*:ЅM�L�����(m$��I#��^(ОU�ƞ���]b��^�kOW��e�F���;��f,� �� 5o������R���[_��������̋'5�
K�iY�B'��G�(�՘,t�U��7����(�%}�"�[��,�20��Ώe�}E�TQ�x�,��c����mk��
>�@ %�U�HD����0Haz��.{���W:��2� &��r��	�'N�F>ڹw!8�]��
Y�����U-ފo*-���p���|'��h���N�wt,���^��f#{T��s�-*�Vj���|VzxDBB�I�M���6E5\}���h����x�ј��;��=��4@�;D�|��|��ߘOu$NW�l(�@�$d��82au��T�D u�e&�S3����������:,��%���&e�	�e���B�$ǖ�x0ɸ��"�Ovh���Ta���/�-k��:q��d�F8���"���ō���%D��*����2��h܊�Y8�W��Js�Ra���m 'G��ʕ��#K�k�]��&eSz7����W�Ly���T�� ��O�et.)������}�H��Yu�����~�1��(��-Z��c�씬�Q�:�/��1W�nq�+��ߚ��t�M�߮��lލ͚,ht�$H�0�p�r�Y��ٓ�<ë}�0�:������mC7 M=>���\|�&��+�u�+Q7�|�T�b<| ��;!��V�6˫� ���;p��<����2�pH�y/:˯���f� Jr<�v9�&��&d'�!���S������?KG�����lwe�d@p9�Q����S�H��Bc��H�E�.������y�
�w/��H����R�W:z�9�ۗT������id��mQ}?	�_D��E,~�_5�8v�����5h,K^a9~�	�G���<9�u���0Q�ᢚ9�Ȳ��<A�3�p���v0���ډ�+�W���ԭ �
uam�w�Z]�7�	���J���~��*V��E:E��1�ŵX���b)?6����+����f��v�ؐ��	�N�� ,8=�j���PR�m\glM �Gv7��l<r�>�*G9o�����G̀�Y c�Q�ʈ�+<ks�> ��u����p ���{�z 	�A��cL��� �F��D�*g�}��lD��$�ˡ�8�#N���\����}�y����s��s�&��PLEݰ�i�l�G�������qn�l�3���%�F�k�rGR�!����N��c�>=�
��#��<
|��*.����"d��U������lK�w`FeU[�I�6Ch���#����L��|�5��|��@�=�������_��8hG�]tCϪL�m=��C���\��&� �?�6��/�4�8�(� *c6��s#u�N��,�	E�>���ִ�2�'��]�ST�#� Z7a]�x��Sig�D�u}3=�5$7eB�W�$C����|�Fj]Ɍ]Q~��Զ��� ��+�4N*% ع9h�7�-��+$���;�E�`���F�2x���Z�yd��rE�\���`)7ޞOE�r�x���
(�E)t�AL�YBF>2ԯzHM���\+�Hi
��9d?�[/�2�apL�b�����,BL.�W2'�{�Ʋ�&�T��gSQ��1���ᦙ��4�KJ�-�M��PRe���㓓��<-G:���>�ݴ|"��aLv+�2	�qw�C�f��j�#�W�Id��=c���Qz�m<l����t���{3t�mf��ț�BњM���v��s�+hf�V��C�˘躰�s��0�K�"I��.n�5�������œ�j�{q,�j� �q"�����PW�c�h��}++�j.���t�7�٢$�U��+�`&3��:���"w�M4��% C�zd�f ==�ձ'y��۳�%@�69���Dƽ��,d��wӮ_�Hئ��Z`�y��/�2%�Lѻ�2�3�����L[&K���&�Z�%6���,�>j�c{��n�
_)����;�i�.�b�x�>S���7M_��@ޤʺ �k�"r'h��iy���@�N�;-�<� "1�}��|X[B�)�Ъ��.�Z����uԠ�^m��O���l����;���T{��&e�+��#��$$�H��ȅ�to��+o+Թ�]'�G4/?|jń�����e��!^�ݠy�H���JM���O��r��*ݶ]$�)�NmX�M��_�es�OH�������<����?��G�֟'��ΰ_��������z&�0�L2y�S_">im�12���1K�����q�|G9�[�sG	��^8��T%.�D��H����A���X�b�7"�#t Q�S6� ����1�!�G�0�3��J"�Ld�k���U�@1Q9]gڬ���L��6Zᰰ�ABǺn��£�G�����y_m���!���IFB�A���ҭe"�V��k'��[��z����U�������RMYO)�D�^}�z�~��lvpj��I�/
����w�όKP�m}��#���ӋؘΚ���5R�"	��A��Ʌ
D0t�y��o�P����u��o\���e4��]�
�$ޗ:o� �Q��-iLE�� ×f��C������i��`��2CM�E�HX�[�w��6rD|D�)6 �7�T�,���K�]����`�4�(Y�˅�4����=��6b�Fj��	�:��8�W4��]��5�ڦ[p;�!�+�j%գ��="���?yĉ4d�a�<�H��.Hȳ/��F�>���|�EPC|Z�ƹ�5�'���"�D�53����������v�̣dh�=ei��h���� �i���&f�i'nsy��֪���$����5���I0|�i����4��B~��b���-�y²�з8K����(���������<��?}v������m+�ukv��5r��.��k�k�|V5���H�-��m�f�Kq��8�U���r�=��#��ǥ���,��zA��ِ���Uyf+�4h�f��Z�ؤ�Ee]v�ч%���a`�7_����^
��c�R�{��\2FS���C#a��
�2�l���H¾O��v]M�X<ʓ�W�<Q!�?_H��9X�)�H2�cJ��vA��z��<�2F���f�nm���^�M`a��p)�?8@7���XG���e��9Q�{{���_��V3�*7�7<z^8�5��$��B,f_@1��$�E�J�;!��@��e)���Z�b)Ny[=4�g��>�?k�j���b�-v�
�#�#�FF�:��8B>$�.S5����$6�Tmf��3Q��]�v�̼�~c��na4`o�[� �����>!t?F���m�vP?E�l�Ϯ`W@�㣧i��g<�/ˈ-ctB���	h~!�O��M�'4Yܲ����c>�Q��Dvh[&�|ͩ{��\+��;@.,��L�j�T�T;�ex$�,���R�ʒ�������b��س��n�	(���D�A!���],�Q�^���>�yI	ͦc	Le���WH4�ۄ�h�)��a]e��?[�b¶n���jF�U�8��B���i��B��/J�\��}YTZ�Ŭ9�P�|d"�U>jt��E6�>�l��=j�O^2��We����g���`��
���f=�M�@Ư�+:(�%�
���{�W<3�a��2œA���|#�"�@�oKp�?:˄���Z��������;����r��0@����:=���tuYI|�=0��>qv'�ɿ`��%Ѳ�}}�q�a�*���]�&�p*k?r|�V�^��h
�M��?X�Eh!�ՓY|Α;l�A*��9��_��R֮�}�T�&��{���"J�ptp1چ��o~�ák>��X{��:#޸��/��!�[��]Y�	�)'�u0�2��@�{�Cqh<�"�E��TB�ʷ�##6���up�q�o����5Ӳ=�Z�B���ˍ�Α��3ؕ+��:=+��-�f7�t>
9���('p�;̧��W���7Z3(縎��p���Z7�-��{��e޸�]�t<��y�\Z��=
����T3Ѐ�9VdTZ7D��J_��l��l��@�r�����/�/�V
F�l,ڀ �cm��?�>8�z}��@�\%�����a���Y`�&�`l�E�+wd���$�}X9�N��w���}��Z�E�E=,ɇa���l�O��i���F��3�!,V�t�_,�WQ���d��"�u�2�(5���LuZ��[���$�+Y�^ܿ�*k=YΤ���F>B���;"C�È�R�A���n��@������2��,��Z>����Ib�����'p�S�C��8����\h��ov��M�O��3�+�N��j@�f,ב�s3�����a+��u��fg�A ��G_?���"��[ Wc������ů���x��$��#�EϿ6�\����}�Q� h�91��<��|���M^&�u�7��0Y�}gh.)ȗ����k���:x����R��u!�LHp \c�6����I4��C�)Z�b X��֎ڶ.��ۿ��@� g� 5s$�3XEYx�� E5�F�s=��Pg.`Z�4z�󭈳�$#���`�2���h�a_�te(xAIO���+z�5o��L���X��͇Ad��-?_�p텺D���.�gi��H[��wO�s ��.�/���j�I����9� {y���?(5վX�5,�������.Im��������]���֮W���3ߎ�A	#۴J�墙8���Mʆ��+c�Z&�w���JV{�ʞ5d�Å�Q@Z���v��y����g�#�^����Q�vOv'�)؎f]lY��K[�4�W]��-�^��*l�.N�(D
�i�w�}tS��cW�4�i�,��ΥqR��JC1yߘ�w$�� :2P� %=�XY!���Bl�x������Dʃv���1ĭ�_�g�"v�z�0v[ֵ�Z%.F�&w����]��ܮZX$^ϡ�	d�RkR`8Ngs�z�|�.�#�yS�S�׼�2A�B���cTVjDR{a���C[�>΃Ѡ��|��ڗd+�ge�]�L�Ʀ�28�[��[�.z�H�z���/�c��}Đj!���v֮z�z����N�`���s0�?��vt��:��ȯ,#�HscPt�W@���C�ǵW)P�
ekf1�ql�������-*����w"qǑ��ڎ���m!�U���g^[�g�#|O|��W=�2aL�1�.��.������-��8������0H�M8��>��ӛl�����)p B�h�軆0�д�&�y'nC7��Yɗ1���m�inA�imk߆�U���sI:�;�uƧ{��62��/z��:�c�������5�[r��9(޲U�i�l�TtF��fL��6�T=���PO{C�9��+�2�~�U#q���[��i��d����{g;옙��O&�X�=���\5D�i3�R��N/�ط>A�:o����u�^d����s�&;٢����Cz>���J��0nŮ�3i͓Ja&Ya�4p�{(����I�Q�hTUf{�(��j{�Y��������b	��EP.��/��%�jK'բ��)r?�u��ח��U�P���fƾ�D��}�������l4���(R���~f�}X��l�����F���f��FB�k�`����h�2���S���Q��&���t,�l�����4/uF�g��,�h�Ss��'A�dr0��0���7��N']5�y_<k���=$�;V{����z�gxJJ�t�2���G)�;zr1h�4%�)�����qA��l����|E��j�C�i˴h��0�B��Q(� hE��S�h0:�ZXI-��Ѫ3e���Z&Q���A�R9�ELFRȟ�y�.�����5��l=Q�-N����!O���r��Ћul���x�̘4IL-�$X���6t��TVYl�Z��Y+��;9e�&T1��:�a(�1xe�~α�W������JIN�K�TY��v��T!��*��5=�����óأ��y�����,�m��]V��wMK�����?�`3�ca��<�y`<"',���
�M�����S �;�l�|������D���ht.��$�e��ߵ�6�ͬK�(�Mݕw�a���.rqZS���`c��>s�AJ��HZrڶ%�t	��$��7����'��I�{�����*M_P��3�&<�˗2���Ĭ�W�ٝ���Y�L�p����S,�A�>;N�9�����1�C�wƳ���v;%f���gn�g�Ǖ� ��Ǜ:!����M���<�{[z�!��0I���Na
�m�w7.1
�,��a��������}�贒�����P�H��G��o���@�.<�V^�V/� C��8��?Bj����T�Ka�o������*?���"�1�)F�7�����Ha��;}�C��
��P����[��~��;�-��o�����9�+�-��%��p���L0O�דF���)�I��%Dv�q܁@��wQm.,�1�-�j�-���KZkT\�@�e�iD�k5�A~cs[kų5�I�L�D�!�E��`��i8%�B����K<����ɣv0) >
�g�(���m ���hmE�f�+�{��bs��H��6&Tr:��ҝ����������������	N�_r5쭳�óW�����O�1���x��\�Մd"����(,�!w{T�AΠ�pJ�$�g��ȰQg�˻l���������/⢼'�����^�@�J1�z�	:�E3s9�i<m�1ɺ:�BQ�	f�䝅u�_��F3��5d7!+�d��h�T{ҏ{0^��#t�~k
��|IG(}"4ɚ�M�?m�s��ʤ���F�7����s��m4OY4�7/�+͜�(z�L�]Ɲ�O�����p���m;�Z�V�Q�8��ɦ+zP��tA��$>��X��"HBa&=EfػP�'�Xk�#9G��1�
�����g�˒$�*��e�ҝ<�����{���k�v��h�4��ZV��G�
����Z$�Ԉ�zT���Cf���X����Mg}*���DT��CY�AI��	v��c����A��l�4�^���9���7��x���5��q(�^z��+����/D'q rv�`�1����yV`�[�p�WA$ ���d�����?��[�����jn���K�ӊ~�����}3������>�Z	Y����H�Rd/Y\�1�3���H�]�CV�R=ǹz: .��������sv����f=�@�~��ިÖ́�*u��P��/Ͽ;��#^>]U;�I�g�d�gone;K5�?<��r���Hl(��u�k���SD�F*_3m�S����1ۊ�~�g:ח�{���^ON�{R7 �)~�:ʹ�
��P1�u�q�>�7�Eu��b��Z�7\������~��u{Yehn"����p�%b�p���ʱV��.6�
�N��!a��Y�lY�4�A��.bU*(y�|L�gS/��٧Ե
��Pա9Q ��83_y��	��%\�Tء1�#���[ߞtʊ�M[�%�
P��s��O�z���~10������G���Ͷ$'��{lJ5�bɽG[Є�����^_;9g���=2te~#��8�\R�q@���@�����K�:C�ҭ+���&��O�ujk T�#۴��䈅Rp~�j��� +ƃr���������3���ۅd�� x:����ke�S�d��Ja(u��(I�*������_��Rwūra��o�!�3���PL�T���_J�S�	@����m���|���J�Z��
�ʥ`�P��|G|��]��@�o��z������$t�*��Y5Z*>\/��,#��V�@|�xyy�\1�)�i6?���!d�=GޏaЈ8�ug�t�d��@޳��_� 	�Ca�(����������M�*�t|��6���E(�h�B��k�\r�D �H�:�6��c`L48[�?�Y�l�kȣl�z)��̵�Qpc��@n�ſ;f+ 2���Ƥ���bD�b�����2̓�?�s`A��ڷ?�i����gX���*�0s�n S8�:n3��	�Z��n:@�l��R���[If;_���|it݉9�	9f#�}-ފh��u�����j��~�d�0���"��y�+���&�6�Pi�*lB�T@<Ͳ����*=!���E�"�� �	ኻԐ��OO�poH l��k=}�@���è�V����?���"b�!.�_+\LO�y��OK/@��&�Ц����/��v4�������	�in�<�N�gЭ ���fʰ���� ���c}{�mA�����TƔ�]!��nqE`��)��|!���qw�s�H����9�X�D��HM$��H�2tK:���s�q�}Um�LI�Bc<�0����Kv����6�m�u�B9k��˓)E�q���c�l�u{�%y��Z�"��oO^�]��0�Ѩx�^��+����ةz���vQ<�F���F�\dnW�ڈc�o@i�y���,C�|�	�W��Vp� 

�W�ͥ����]/�9�[ó��ft@i��f�mI"8>�kn�� ��c��*�A�vuQU���]�SS?\��^c����w�A$ Qz�}w�{���~=��k@Gau�K�Q��!+���}������]�azc��*����@8�XdԴ΂|�&��w���69>n�0?.r�D��Bc�a�2�L�nW��� �s��3i	��d�\*v;��+:�� P�T����i��	M�Rd�a�D%���!�2�CxS�3[�Lx���\�t�K��Qm`a0�� �1��'�w6aL��D˴��c
���[�Z�r�$j���㘣��DIѐ�s��87��!���:�7���Z��JG�Aq/�ʠD�;�?�&mx>�c���t�美��4Q���(���a3�+�H�=v	�eT`�3K�oh����a�"j� _�K�[�9�y����S��٧�.����P��{���HW����� ub�(���tf?����#��a���"���gְ+������&2�KM�~�A�ٳeq���ƦX�00i���a$���7�4�I_�����B�}���O	��q�ŗ5���'��"Ln�Z��[0��
�>w����=���}�_.�6�LL�����=���=�>�9izڜ����\宵i��w����I�{�|�H�"�*��1e�l��[!&Pṉ����f�ɷVs����C_���S/������{���5w���" #�$�v��.u#�MK�B�v�<�h�za��;k�G�ڇ�G.��걣�ud/���_.
� ���LyO��)�B5��[�jT?�p��T�v����)�u��8�"Z���5sVm(��/6
�ls�z��怶I?k���Y�jf�l�ǈO~�h�/Yu�iq��87�8JxF�\���B<���	(IJ&� ���XI��'U��?��X�^����19Î���-��މ�偧��ᩍ���>;9�j��P.������i��m�r�g��s!���p�{�M�^��T�� �"����~ �QH����suR��)�9�:����V��L��=�L���.P	�0V��7����ķN2�9~�$��L���\�`�Rs<�����'���P8!�c-�:hl��_�x�>[��y6��K���m$5ixn�=����;�Y���?	�N���e�f��p�ۑ�h�fcx1����!�D6�C�X[>k�u�w-i|��Z�TQ���}��_M�ݵ1j".]��ι��N[�u�B�qPx�:um��>���ϔ������0r7���t@���`�	��J�����������y	��x�޴R��#�������_kq��v�f�{�i]��v��m��P�	���њ�b�W�	� ���\�5��S���ǘ:��2�'�L�Z�$�ɢ@~4䶚x�V��,I���o� ��?l�M�t{�eĔ���w��X1�9o"�'�*n�ೞ��7en+���L��`;�V�pX0�2Hf��ʭ*����~����8�W�q�ؐ[,�e)m���$�𡚥{����,�x�\��|�M�k�>����I��3�
�\1'd�T-�Ƃ�w�r7Z#?Mvh'+`��t(���m�� ���FS�hO)`Lk��l�4V��b�d#��-?E��L�3&L��9�����5]{�GC�IY��B���v����D��M�4��V3��
�3����HH�h��_�x�0(?]����3��ub>o�J��9�XK<<o�Rñf�V�q{�&�"*;)�b'���1��&��~���ۏ����l�\�S�������=�&��Z����:�_�i}z?14�^���ܨ�6��"`�nM��"Q;�|*�l͆��\"�Z���M%,1~QN�@.�+a#��)�Mw8Ąkr��n�.���o�ލ?�`Y��
M,N�ҍ�����mp��:�&�?ʽ@���0�Z=���Zk/C?�WcK�b����>]7������ �kK ���ʯ?��[oڊY�Ld�ju��w����eu��rm )�\>2��BZ� �"ت	��Gw8����g���`	+�?ƻ�:�9�-j�gs�d��6����=k��)jjqfsb�ֵ��~+�^�+Ю��D<��1���y-�F�<��BBx��k��N�e2����b?r.&e�.��q����g�#�SF}�11���������퍀���}��V�����Ub��E�\3b�c>Q�L�#�f�%ا�S����:Al5�
e:�Wk�7��ʾr|��pL��{"L��wJ�w>X,�G|=&,X���c2E�g}|��+��X���-����l�{|B��ίl�����B\��+�%����M2�`=DW5���p��H^N��������*w���&�!5�������|��4O)�J�
ܯ�<:��}�� vL2\Lo�&�H!��0 ����YC��ĵ1�#��$��pF���G����K�+
3击Xv�
�e�9D<�XݪBMN"�Z�j��EG�>iEx�2\�����D����LB�O��_���y���Ӆu��	�h��hv��B��1�����m�^��E��I�;Ӵ�
�Q�zǭ/59)/�w��eL9d\���R�|����?{��!�S;?�{3P	s#�/�����DIō�w8z��Nq� �S�RO=�#��k)*#�D�f+J|���w@0�`�����8��Z*��Gru��2j����XpźCmLz$�Ʉُ�{V%H��`����_���?�����f�������lIh\`�}O�b���.�w�S}2�*�z���uv���d���3���	�mR�G�V��&y<�r�8 ܭOsc`�}���-���(DQ|����h�49{�z&z�=`c�7��(^h ��� -U�����e
�r�� �*�3
���e�}FR�x`��O8�#z��Ѥ�_�j��֊t~^��m����;�etr&�i��J�����KZخ*ce����V��)S{㒆�~�/a1�9�>�R{��A3���cߩL�ӳH���7�h�qp@+^e`G]`53u)�c�j��vC�ӹ��u|��by��m� q�s���g�n��M��|�A����}��)J�#�����|��������\���l���>��Cz���tA�X���W�5*���kd�)�����,�o|��h�]��'\02]���4NT$����.<�qb������}F�,�"�@�X���Rr9��r�hHX�%}�>=u�)Yv<hR�ӳᓢ�ə��#��5��Hf�ܷOe���8��qxt'X��^C����?��L�Q^�ov$�Pcε���I �\�F����ͮ��M��z����j��٢�ļR�u9��H��f��y2-438���˦&�yֳ����pI�V����Ͳ	!}��)ȫJ{�KzJ�#W�b��[���M��3W9Dv�lśu��%��[�]sc�4��r+��Ra��1�����4(��t��2� �&%���\a������QLf��MI/�R�=bk�K�S6e|+�]��i���}��]�=��w}Թ.�l;/�o:�JJk#���
}g#�J�|1^Ƒ�V�}��,��p�v�*xżHc�*v�	�$dnnѣ�h�5��ӊ���	������gm��1>y(;~HS�C$�����!vj��i�[���v�WR2�)t��,k"�fCvݎOR������h$j�%�zUw�G���G,Q�6iԃtH(��9��T��/��ơ�B��W�����3đ�^��$ϳ��TJp=9^$\����Č�b��ث��j�*��,[�i���H~��ꟾ�	D +_�+��6�R6�φ̶ɜ�
������P���c|;!I �I�r���d���"ҍ�bQ���U6���?��A�B�q�_�Y^��'!�
H�H�k���0շ�P6�7��"�Ę��PE)��ܞ�п�?��?]�^����L� �a)�֓.�؎�*��%,������#ڽC0�)��%�Z����[��ʤY�ꟻsp���,�\�4֌��Tn���� p�Ѡ���o:6+�ǜ `��Z�/��R�[��~oʫ�����~�t6|5�����(�[��Ig,f�~S�Ӏ�
k���Վ���W%>I�=�-��v�W��O�'�y(�s���*'P�ѫ\�ه�Ȅ���\�Y���
��RiOX��\�R�ɒo��e������H���}��;�i�J��R��;V��6���f�b汿c����v�\m��v�G)E\���5�3�d���"�tW,�K]���ZB�E��0�g�#.�O]��B?9+Ox�pBx��ͅ`��&��߭&=�F-���}c�C�N�b,Qw��a��n����^w�q��r�w�xߝc�6��c��z��'�����@��&��t?�%8Y���8BG�z},g^�F��&�Ű��	�E�0�G� �(#�v]�:���D��ѥ�Ry�����.j\aa����1�U�m�$�fܔJ�ۙ�	��[��t�+8h~� �;�[��9�*]����-Kkz��51��+5�qE�ט�Ymv���u�)75Q9��6{Db�J}�kl��G�g�3^̤�Gߟ�G��Ғ���_�>GU4���g�M4R��G�ߥ�ɼ�7�����t>�S=�;zSP��j�f��g;oǑ� ����=hO��d��Ln�[�2��br�)�I�	_c�/�x����xwKH���}�P���dY�����#-��܋)��T���u�K��u�vt�Rx�q�r���ʤ�[Z�'���c&���BDJ>mF��Q�i�:x�t�Ϯd#a�gr8c�`Tx �	��9Dp�4��5i��z<3 F3{(k����Aȁ���(R��	R_���oV��D�xr[�aF������'_��ἴ��=a�"�!p���G�MP�Z�>��C5>Tr�-�W c��SHo&�8	9�F�7[�y���?���tgx��Q6��M�m�^r�%�@Rb���	�f��$[��r2˔Ɓ�:EVش̲6��|��X��#B�7����������4�0�OցYIe�/-��D��+x�t��*3,�3��?������u ��!H�48Ь��.�zT������=�t�����,RCaQ��lJ�tP!Ŧ4��F@��� ��'8�S�B��j���wi���k�賬�G�p��h���e5�|}@������}�b�r��f����P���l
�Pp~4[M��z�hw*�+I��-���� �ȧ�4��o�!	�{���;07,��x8�x��D�B� ���$��ٖ�g�N�,,��e�T�����.������P�2m�����n}&�n���@9�>� �0�ʌl6��9"����O,.�����K	R�\�9fb��2�<��zC����{I�h�z{���,�A������d���߀��H�y���!������R��H/NJ��>tL�tݳ�������Ie��_O ���׃h����H2��uC���b EI�j��&u6�����gp�<8�s�l��s���bmϬQ !�HТ�(��)�i��.��M����+�|NK�S'Љހ94-`�$��\����*ZH1��[�,s	c�U�h�k�PɈ�>1Ij.���_ �~~��dM�[����I�e�7����ur�Q�܇ѹ���*�Q�Q
�z�H쁋������	 �{S`�p3aG^��VU��Q��v�;~�A��Q��DG1��Ą	S�@�����ʨ�f����Ԃҋ'g!:'wG	a*���v�nS�(�3��J7ed����>���fb�p��O�^7���{��⋻}&>��:j,Ww=6��-5��b���:nW���b`��+D7�Pu[y�T�1|���Ѐ�v8��־���L?�r�-����&,�`*05�e�2�i���w�`���w� �������q�Vt��{˺��n��X��xF����$�I�l���,<V؄�W ��r��oɩJ�7�8���"��D���f��մG|�p��i��]t�J����W��%��4�0��iX��$���λG�Ͷ�&x p#�Yߤ��T�B�@�"��J�����Z�;�$a4}7l�v�V�d� �ˆ�� �����y��O%�I������K{/�X���on>$�w;w2D�	U"�;3���u�v��$��͚P�w{��G��
d{�)��=�׳vh�쯶9�����v(���'��R�>i�E�� iZ~劖��Ī���"�wxj����X���jθ?M=�6���&LeH�i#�P�l�F���a�����O�#�������#0��BN��,�����mX��5	;uF�g��j{�*h��	m`�3-o<r�?:�>+�����2�a/�:¶�{�rQi/���F���� u��M_�e>�oo0|(�i�^�J���7a��&3n�3�z����/,5:C�%.�kŀ�g��z��X�W�`̞
9��T�5���@y�1Ut&��#�4�"5j������n����:�X�l�8Aּ��;�6��5�83M�����6�X��SU���<O� �#'㴴6��"��[�Zs��!�PZ�3��bo1� ;W�*��}��Q+��#���H�!)?cȼ_�JM�����gt�LKW��U���l��i�L�L���1=yȧ�,x9��[F�}��1}�Ūon"��5V�pፔbBE;����!e��e�#��v��d����j�����O*� >�>�0�;�����۫�#c^�W�B2[��C5v���<�������$��+1H#%����%�B��ߨ�^`�r	O���"���P<�J��I�X�/ͮ�ȫ���M�Ȝ��������zu����ઃ~\�
 ��	��y�G%Ⱦ��?�ʼ��M��
�F�؛�6@��_ƾ���H�$d��gm&%�w��BPN�s�޵ a\Z�3Sm}����RPnPs5�mb���^"�-�ʼ���ݷ�.�֋��Y-Pō���a��
Hhو�>V0ںq�^�������Z?�L��F3�F�r帆�L���dÂ�q��GJuḰ�'�ځ���q�G�5��ӓR'�O���4"6|�'������Ň���궨�K�!��2�v�V\us���0��򹺴,f��?3���u�hR����Į�j���PF���e��%��h�̞@"0��8qML�9?lf�)*�c�9ig��(极^]Ԍ��"֑K���$�2¯�E����wEa)��r��?������e�˸�)�e���Ǎ]�
�+On�_s��b������_G�}�KhB9������!��K�ښ�@_�J�h$�M��A߹�C���LUg!c�(*�v	��o������E�fe�Y3��\�.�u�g��u*E�X{9�P�t�י�l,�h���p]d�i4cR�搮<4ϑ�AE��3'}�O�G�BADc%�9w�9����V2*˿'T]^=P\�L�X.81f��VNA5/,U~���f�&'����o�{��F�K������K�g� !8�O��ކC2æ�b����*%��~�>h���l��B=*P&;1jƬp�88���s��#��k3L_�c1�n!�sޣ�X�=���.�l����ǇF_��������f:J�.�攞è�tp�\�v{dL��]�{-~#v1�D���h�;��zB`zo��6�U	���@p�9�]�/@���l�D�����i�^�5F"��fѦ�f.��
B��"@a�;����a$�����%��Գ)����y��2ՠ���p:tI��3Ƭj��{R�A�Z��C���9����44l(�*��G��=u�҇S�Ḃ�?�+����
l�k��/��!
���Iڸ}�x�������Yq���9J���#y�s�Q58�:(�Y���e����#<��*���&ӵ�����J���-��L(�DS�������%�b�M�@��i�4�[�)�+c�{~��@PH�`NU���dOhsa�@oL=|�� ɓ��*�k5�$������nNr�MqL�Pb��\�A/�J�������tp�j���Gſg�O��V�D�5	�O�Bռ�섦��-��d6Hs���;�w�!��:&�����Xn�婏?�XB�.=�JTV��L�d�Q.`��aOUb�MHI�xdeL�O)<(�v��V���T=t� s^M�k��}F��\���	x��i�L������܈�
�\N��XU�$4˩�%k7��{6eB��`Z�NĊ5�JUt[��df6W�rh"ͷ��	��2�˂>
a�
�X��7����V������i�d���X��vzW�9^n�ܖ�.%c��>v�9�۪'Y�©�Rn��b�;�|���h�L�95�I���1�;�B���M�d�`�e*-&�[�ʞP`�%AI�3G�e4��� �O��`܅�"W[���|�z���������;B���p�x����0�E_�Q_o�&#o�w��ͭ�ta��el�638�I~��4����jt���f�% #�=k��zlA����4�Q�h&�W�� ]%Zܒ�[�Wl U��2,#�A�/�6=����ӮY)֏mU)K(b�s^z#{P�`�����d�
�	��4�lb$w�'����˝��됹>>�UL�>\j$ י�l.����"���Y�J��
e42����(I�>�*J�>M).�
��YmNV��%;&-�Nؼ���R��|���5����ѵ����R�����M����<�?�3�=�b�����g���7�M�*�vBI�N� �Ѿ�S�������!S0�
���M'��Vx�{ tW9�\!�Nݿ+�l̹ܪ'���Y�]]�Z�@��_S�b��,\�_p��w	㲞��R̰x�^�����ԝ�����1*�LKH޸!����S��/] W��t�5�Q�9am�������>�I<�u��\i�b�y�\W]�~�߿[��L���Zf��8�z]��!��#s$4�3�=�#p���}��y�hH�%+���k�vX�+3!)םO�Y����,ҋ�1K�H��G��>]���ٽH�_��/ԇ�� &K.�T���	A ����/KD��8���vĻ��/����(�:��|����J-�4W�ȓl�{��~`CN�F&�Pq�S���;�����xJR�<���l�U0[��H��E|	���J��6��"�:(�gٯ|ot�1a��!�ޒ2��mj�����vp�8�h�Iꚫ��1�9^��&p���z�gR��Z�M��7���^�K@f�q��ʯ8=�7.�i7��J��'�#:��Or�,�2�
��_z2Y��8G�>�a��䩾y����N-M4~S�Wم:��X8�N�Y,RL�~�\8 A������d.ec�x�j��BԢ����B�-��Bv��Z�ׇ.;F�"Oώ�A�\"}G�1��I�}�T��Q�����kW,�&�P��C�F�+���ǎ1<R��> �k�.2�?���On�GNK��u^����طY�囸�"
{�O|Cf�	�E.�����`=�\I�S�:�W�k5�藷::|� 1��tIB���$F���!Y���~�G��*T��Þ�N��l5t�ҧ�"ε���N�s��q
+���d/͎���o���x)�s$��o�@�-SIB�Ĳl|~�Q��;3��Rr�QU����}K���9���"�o<��H��f�=�U��'��M��~Ik�� KW��J�Cp+�a��k8i����}�W�q�����V�D�ݦW;&T]�y�����j�	@;�F x�l�wJ����p��&m�=KH�꛲C7a �h���6}�D�!?�ν��>�GK��7c�(���؆�e��xG�����N��M�+���VI�zj��b��Z�own�B�
6��tɺ8؜SrCu��?��9@ vA����Œ�5>���v�,�Ajm�r����X��*\�Ge� ���f�iI��'p��@��0��{U k�`��$�m�o����M�a#��B�|�]�(t8�+ŭ���G%�6�~Rj9z\etI�$o"&z��{	6�� ���D7l�?I���T�~V�:ȩ��}��BX}z��"(p`D��
�%�2_� ��ڱ��Ϛկ���c��y\O�P�mGS;`���Fq2
�� qud7^P�}�{��O�7�:�_��#{�~O�?�{�>g���1�k�A�����q�;-7�C>x��"KF'|�Iy�s��?5�r?�ALDܾR�[E�m{Tz���1�`�U{�{/���ti�xb�w�J�/P���o�w�Z���f��1^H�� ������V��y�~؜ejb����OC�U�6�IXa�m���R(V��CO�� 	��򙚠��g��R����.�����1z��/�������畺=C
���Ե�?