��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pd�Ύ���yya�[53㿅`�@�r���m��6��n�GW/w���Y��v��z�`����L�2'��ցy���3�{>��Ŋ)LQ �'��nX\
`xʈ=���q4��b�3�[ĭP���S�x�l�0_�>�:5��r뽳�8n8�^��}9헹|�K{�-���`��c�Ȅ�	~�q%O���A��� h�3y矰И���%;Hqj�_�+��꿾hz�dG�M��})=��nsB
�:�ZJ0�2B��4��޴�T)�o:���g�w|�N��H�''}=~&7W�؅yT5);|��e�(c|m��J��H�����vy���o�"m(�ޚN3^�ȕ�Ŧ��r%��'s��T?��,�b{�|�����N�H���:9\=�:�T-A��FZ��{��,O�/��S]b&XY:����S0�<m$I3ҟa�1��M>R��@�5űM�7�2���^���
���aa`�coyH4���I�u�_����l��L���>ɮu��k��_|>�U,�̰���1�	M�9�\>D��a;���2�y	h��ۍ;��PQs�@���éc�}�\k��F�|\�i����#�©w%�Y��|O�m=�K[�wi�g1KW�ڱ;#���k�"�F�B1gR�Ρ�_bi�:pti�V¶I��F���ԧ���A=���DXﱂ�y ����+�v���8㫙��c��1��K�_�������3�Q}Î4/]a���x�G����pn�v.����.WV�!4Q��е{���A��|� U?�� ��洍9R�����隠 ��G��������ϟ�u!3�d�󼔻�a��Y���ho�����7ݛpQ.�k\s���|�K͹/��4f7��a�K�/��scS"UyUt�Ct����`�i�|�oل�!����W;)�B�*�:�
w街� ����]_Yuz�ulfb�j���S�k�ǙT%7���IC+��H�gl�+�K�bE'Ws��$@Z�<��<]2�=��ކb_c����Ϙ�\�?��,�����������(��"��=L:q=6bL'!9���q�Di4W����E�yL����%�i�k���Qhӣ��� �rmD�����\������ɀc殉J����1=J5��o����=��!��{���%�Q�s�� U���-��0�eI֮��H�=�q�j8E1��~z��^Y�uի�e�����~�r�;�l����
M��O�.�^��"[܊9V��s��h�1����������\	�
vV'���]�'��Э
Zґ�Bq�9���a���P��q3���u�U�|� ���c\�O>F��w��T�����'�J[�����i@�N��Y��.��h��b�{0?�Ң��?E��@�Ʈ�i�p��U\M��z��9:�6u\�g�f	�0ZCV�����"�꾰��>>�\��a�9,繟��-�  C;+���lc?����kw�:� dh�6��VC������������81�n�d��a�x��^P%�3�Z*oz�}�eb�00 ��qGANR�����NV[T@P�M�w�s��
�G.���g�N��'4�o4���Uϒ�g"5q�7Ke��q]J����*�=N��q��/޳���"!��W>�.���V��
�V��f�`/� of���w����nI.N����I��NO�Y9\7h�%G�C�(�� �g?���k��`]��L�@�A�M����ZM�\�OZ5y����]X�ނ��l V��t���e��.0^�	�y^4M����ɽ�a)m�vg��WE6h�v�X�p��\�-g�;�\���Ȣ��H�&/3�'����K�c��{�v���j�3�)U�E	�~����
V���E��9���G��0[����lV8Q���Ej~����P�ԣA?��'��M���s�E�vCqK�u�Z�AkǮ-
q���h�2a�I-��˂pY����qq�C���]��9�'/��R؅�l���SH�ݺ�Y �#)�R`ޫ�y^���Y4̺�Ț� �^�t�}yQ����3b)U��
?7aB=�V�J�2Uv�p����h��\L�z��� 1�C�G���e�
}f�֛�����f?m^D`ۮ��D�V�b�Y�oo�61�}�x��r��S�g�*[�ӯ�� ��,2���3��eu /6��ĺJ�0�J�ա�"�O*���%P���.fZ�����ԦH�cw�@�zģ	���MϦs|�'��\�j2�C���y�Mm���v�e< �	I�90)a���{����i0��ќN�@��|�F�I�m�H�2�u�� �.7A��ͱ�w1E~V� Ϊ�4��������Y�N���7@����J.�?�ȅ9S��"�R�	�
8�=	@���y3V���HM��*�2�\)�=���[����n�q��׊S8D#/߷dM��	�l�OΩP�+I�kʃ�!��e��f��/]��΀�M忻*hak��ˋ-+�.7�ܗF|2���i��DFIXrk�Ch��H��;�n:�*J� �>]+-�U���_zxoj���+Fg�d�	1�/�!C�E���JtB"����@fr=#iMT�>���n��ݑdW���+�כ�]��<(\`SA����>� ��oqp�.U��J��@kTWV���2%��b�ۈ���uOtV:���g�з�tD]%(u����ĢW��i����?^��nR!N�/��=�x|�b�^W�.�%)�����8��G�ȋW���������9�c���w�ѻ<��[�+���j����RE����=�4��2iM��<�K���m#����p�D��s���;��y�f,�C��B�nm (������Y�:�ov.�$n�AK�N��n�E��@��s\�l��4��������=�����P�4,�AXe%��{+0��4�d�d������̋|����fpߐ>晬C��6������G:�����ڴ��6�q��t���G�煁��SP��w�*o�mۣ��ޥ5/9��k��b]=J����L�c�B�@r(�깩P���˸F�|Ff���&�����G��c�0�͕ϥ��o�F��x����Om�Kx�L��w�bV��~��t7`��AJ�+���^wp�c�w�Q��5���ǈ��3�7���7Ef92�]��Yv���m��땫��Q<F������A�m���8r��7_�����$㯄��/
A�ei��~�`�[����lt���V%^u��Q�\ؙ'��N�x�{zda��Ue��b򃾥�g_tDq�'��-��4VS62����݋ĂbM�U{&�V]��MڣX�-J[��%����S��ρ�qV�w�����#H�л�6�U�!�����h=��P�%r�߁3u��R���Y7 gQ�����U�+y��ss-��4���5R=x�$�6��6Pm�w~��LJk����� ��,�����������-]���=B�j�u�y�� 
'�\ٺX�u�}�(KY����`���n��	mF}��k���_Ϸ�wR�E�h�(
�Dh���d���jv��G��SC�X�T�X�������fFf��l�L���r�u�kM���r���%��a����ʢK�z�1��x�I<���ɱ��h8f�ǩ��sZ�E��̵��ƈ��n���3�k�;�SHQ����h0�uK׎��a��u/�؂8�J���:|qus��� �eO�uQ�UQ��}���t��Ţ�T��6��C��׻�i��LF�D̫n��S^i���o ��h���CDa!���N�� !���ɼ4ȶˉT_��@?�����|F1!WP��I1�?�2Y6���+������������u���T�_JƁcǰ>�}�뢺7G�A`_|���G�G�Ɋ�r�ꃜ�5RnD���/��@Ģ�,<SWnW��ķ�ؕwJZXc�eK5é����x��v�^m���l�69��(�R/�'q=��'S,�(��~=b����
s�p��:�b����j?IC�F���I[�(N�BS.F��e�I��N��=m�{�o��LO��7I���;�;�ں�嚅�d,���� ��iO�-��L�}!��<��(���s�ȅ�1u�**j���M[?���:�Hʍ"�����b3�(�уZ]�Q�w4��[ﰔ��z�gx"��C֯�L-���R�BF�+�T�.P4���&&���`��.�ydEM?�c�Isy�v���/y�7����6.���lp�Z����?f���> �h�H7�5��L_�r�1�~Í��5����F��[O�z�33����+��KpBe;n}�Xil��$�'R�P���W|hG��{VW<��K�ve����ہ�zը�K|�bV�fr�4�J6R��(V�x�zJ������A��c(^AS��!g��PN�W��xa�/L���1�Ӛ|ͺJb�ɘ�	�?�7��vȉ��K���-�<�>v���J9x���������0�u���`�U�zant�\٬��c�6�PɢM�4Q��s:)'�â)�O����#؀Z�,^�<���$�Ԡw�r[�}+�4���yF"���7m*�k2�K�+�=,J綾���M)\�j�����[qd�&��#(h ��`Q�+d�en�5{�`m'�em��C$j��&�f���3|��~ga8%@��@��GYۛ��;�g�r�79��=��)Ք�`0I�y�]|��iy����9�O�瓹��w�%*�?
ǿG�d�{էӾDh�b�#Á���]��[�cϳ5�}�mE�%�j����93o��*z2dx���Ey�J��(����;�D��o!@�� ��T�M49jR|��a	�y�R�9b��F�켌�z�rx��F��|���B{E��rŽ�՜:%ۺs�I5#�1��Ҿ�$,�s�To8=_#xM��ăH �A�ֆ�"�����H��=B��:&�}�0����Ͷ�0e�q�a�y h2��	 �	f�:���'�7ud�,�y��*��6�ەb��!^�t3$�/Ow�?lX�9ۅ��	�լ��Z�}~������&�0���_�["[��F� l�`L�p=�O�iس��K�q_�1��%7��.�������jiXQR��LBf�r<�Z�%+� ~a_ǀW�,b�8|�߀�3w/Uq&93���5��s�UY<1�"���|��b6�_(1>4(��+ �����}^a�+��l1A�~�U�_�h���V��[�F%�x��W�S2�
n'R@�)��S*<��.xt��Z��I�K�g�%�9h���V�`w#�x(3ʗoq��0+�[��,M�&`�ex�?��2����a3�<ۚ(t����2F����9�ٯs|Hř�����* ���~ ��1�dD,�m.C�S�C>?/)�i�4����+����2�����F%a��{TK�z�s@��D��e���{/������FϑTZ!V/O�Y�+k�82E�4��x�2ٟ{e�Y%���J�i5��X˫l!�t�ZZv�b��l&+V����1��f��+��Ň�w�+�į*�%��^�&�ƈ��9g;:��7WT#��=�#V2daɖ�%�����f�/�h;�g�'Z+'���j9�����!�d���j�-<�$�Q�W1_��+Y��)Sr�BrqnƓ3.3BٷM;�S��A��x�bK���H3yg;<�����j!�nD޻���v��Z��x�)'���2�ł���]�a��6�%4���m����4�ÝFɆ@���D:�U���ӗ"*�v�~�\]�MĞ��|�tϖ�@��C+*f# ���0��ٿZ��75\ǩ�'a���hV�bM7���,AД9:sUuzS �����of
{ ��(2��V+���mX��e�����C�~8��u�TA5]��[~�VWy7�8|���h:��1��^Mg��#i�\�\��i9����V��z�՜#��C�L�pU���;��F!� ��ßmc���C�PD�u!�0ˡ~�ܳ	�}=�\@�}'�#����i�Jif4�J�~!�"
�g��-CI�|�޵�[�\����Ȭ�帤�I{> n�mM��M����()v���zg�84	�S��6������ |�Lt�����J�#��O��9����ĭ?�p���&���W�U��pab�p��6h#�j4�Q?�j���[9�X&sy�d��5n�*�~���3�X�ҳ�-<:s����j�X) �m��^���K� =�w�< 	;���.T6~(�ơիV=��¶�U���$�H�R9��Y�	f�NA��-�t��YoeP#ql��ʢ`�\��N�5�8?D'C�"�5�L��5���=I�Y��)�q��5d���Y6�w������ΐ���
��|�T�gޥ���O0�}�� M���#icg��{i4ű=���8L�cs9���_���*Cy1�hP��P�:k���![��t=	�n��Ƃ-f��~��'�]K�s�i�	L�����W�f,���n�fpP��.E
��vc�P��Qr���s[ۑc���rfň(P�I?���G��ܺ��x	��a�*�fݬW�����@��!,��0 ��F-�7�F����>�l�i�s�3ņ6�~��P����ʏ��pՋo�&�T�\�a�ծ��<�I�`���_���QzZ�4���ʏ�:��(){0+��b^��U�qy6�)�Җ�p�ӧ�Rl{���r�����r#~�Yסh>i����� �n�2h�+*�Xm]r-���&�/r\�ё.�v���^���C&ڼP�}
���{���!�d~�e�uޗV���*�%g~�D����2j����
�-���Y������֒�k�'��]�-��:�Yy�K�v8�:�]��>!����[�3�Q�7�깘��^e�)��l�B��Q���u�&��.���F RU�Ӂ�$,.M�ZD��Y�`�}͋��`"�lQ�v $�?IV������^�f���)��?F�~R�I�*��k��qj�df(�w����q�29-�k&�IH���t�9�x���4$����~��N'wEO��ƙ���ڽ���4�ZP3��`t����gFT�X�>������8_��?�[�ebXt`c��x�W�팫�%J�:���	c�n��-��w'�pR���+"0O���k��o,���+|��m��)�������|�E"|���0�$j4ṓ?a���aHi���������O �2�N0XA]�.`�:1��g:ɷ�u>M	��D
�]���c�Af9�=��	��{���u)�|�E2sb�|B�`6�>�!����NA0�l�d���	9���]��U�z��n����}�+1 Ho��W�ٗ�-�ִR���F(�����ׂ��A֝H�+�>��zTo�ϧ}(���+m���:=�˦�.������K�u�h}��B�t C���7����k�~���enzt�h�*�DH�Jp�k!B@=���ƜAaܓ+�"QH�Tp1��Rm���1}1l��}�[�[{��O�,��m}[O�dz�+�?�$�R�e=�Y�*�n�p�n��Ď�0�篫h:L9֧#8q4A�O�z�d���5�zG� �a-Jnk���qW���G	�����dX�dK��v�Ag�;�B�V�R7���rB�ޖ !6�q�l��x	 SrMAo�Bv�CHS86}���~gV��?�n;��E<�����υ�ie<6{��J*��y��������(b�v�%��\|����Ho�1�������%/8�[�z�1}�M�=�����ǔ!�w�jx�ba�g���?��\ϸOA���VN���Ԛ�%I�I��>˟��9�#�f	X�� ��8����W?�(�:����j�����#	���-n�	�(�����'� �G�U�S/�t��'��������P>�lRɱ�鑅xH������A%�boC��_Q5��U}�������o�N�O�/ὓ�}�����>g[�Cb�Ũ�h�D�|O%��E�?2�u�]��&��)�j��E}��=�����B��K��a��G�]�W]]���������E>5�(���æ*i��vT��ԑc-�^~v]T��5��I�c^����)���V9���;�M9G���Qu�>�$	ځc&Y���.2;��7,;�9��.��[�J������*�F�F����Ts	�G���;�ۊ1[��q5�oD�}l��1X�V��O�А�8d����o�?L���jY�?�H	�_���]���/]&s��̚�	��r��f]��A��|��kg���<;J�1��
�f�˺n^{z��T�r$����5�oh���w� *襆 45���mI�Ϊ�@�
cq�`&��+�>��#��|r����]�j?ԑ�<1h��WMlj��q�t*�!nP2сL�uA���wW\$/��r�E��6h�X����dEb����G��9��>x��@�Wyg�Ϊ\��;�IUt�z50��:�R�	��M#;���
E�G]��RC��=i��?�4u^��\J��o̸�K�;�����}�*��j���t��IA�n���0�����<�XB�[7E����9�?锵��;D
����^�]#,��B �mmEL�_r�l�S������7���^c2Ҫ@�S >uY���9�i�^8�8FGd:�㪃G�[�^| �3�<�J8�<*��2SϏd�07��8��1��O)yh��
�tB�`���n N�qŨ6�M &a�J[�c�̜c�J[e�XG�IV[���)��C?o=��݋OJYJ��W��:�M��E#|�uI-�T:w"aI��=>o8��흎��J'���S�㧁.��=���©|VV��A�yq^�^�d��*�{��m�0Ȁ�ŏ���3�+�Vb���f�OI��+��ʫ��!W*�L�Ŕ��%�Z���G4�Ed����7���>��ۢ�P4�T۞9�h
vv��WL����H\N� EN�7�V_�
��������E{�C�'j �^��!Z��`Rvŷ.'ߚp5c<�<Bk�ϝ��׼
�9�� ���D�����|@�����f7e���Ruz`bJ��D��m��/���]�6�G�T�A=�풇G��ƾ� �ԯ/vv8�
���ݕҴ���,[��p��wp)�����S�\��Z�6vw~JTK﬈Q���A��uI+�?�|<.��B���88�o�Aj8���l؜��R8R��,�䖄
͸����\r�2XȢ��c�<Ԛ��N9�����ѱ�TfONf	A(�E��6>��b�|��t&C���#��5�� ,�=��/���$3ξ��<�xd�J�� G Qy2-��G���!�N��PM �F3].r��0�5���i�i�HDD�bC�z�ҥ�J��ܱ��|�AZ��ޓ1xʖNa�a2ȥ��$ՠ�ߕR����)Oݱ���$���.�l�ֆ~2vl���`����&q�U4��)<�}���N�������+�^�T%���M!y6��@�p�q���2T�? �b��|�P��r*A�@<�lGa38�]i�if�`d�I����bL��^�R�N�U�&>	T���m3ڍ�C�����%���F��0z��a�cv�M���Ͼ��<3���vd��N*4[��h�f?�"�
�|���U�O��&i�����4Zj����W��/�M��E��b���C���m�z�[��c�B�| h������³�1e `�w0�%�H�f���1~��x�xw��vh��o��O!8��D��vE��;�p�3�KE�o�(�T�:V`f��E��rD�!6#3�����@~}3݁�N?�����bEL���r�V�m$)�G��Y��  &a�s,�4��o�q)3���J�'f�P��9ˣ�!Th���̅�.χ�u��_|Pr!׮�,#=�Yh��p��qwj3�`)��Kڻ����I]�F6�*�O�{*��0��)\���R_	�^��]��
w���i�
�9uW���o�,�(��(!�k!�ڴ�6ł���<��v��c����e�M��)���wW�]]:�_6�,��kC���1���ɐ�L�sn�8q)X���8 �q�&^%O��~�o+�g��j{*b�B0�Y4:�a}e@��fca��|�	�u��$'�D�T���o�ϊ;7)[��f����O�M�V����ݑ,;����c�7�U�6��;��}k
Pj�fّ�Ђ��jFg��8`����ۛ �ژ��lA�cc�o�S]
9D��;3n�7��X$uf6�W�<g�V-;�{�>h�^�*�.����OT����R�*?j�R��T-K^��Xh2�vx�s5y���U2'AFYYUŊ٢v����`ku΢e��J5��Ij���+�/o*�Zǋz1Z�jr�Ja���=�¹J�����>���$}3�;���g�_6U\u�8;
��Mt7�f���^0����hs$Jg\��L��BL���7ԛ��e�ΗD������S�sG���7ٗ�_�4[>���l���8?�C�ʢ���ht|%;9����M���wGJ}��#��2#!&���ք��}�I���edo���v.�ȖW�=�B]6g�b�����ο�0g����ÛCt�S~���P*��gK�v�v�k��D�t;�����Ѻg�j�%3n�]�|]g�9d��^|c��T���Ϳ��j��<������g�Īބ���O�1�ᬕa�U�֑{�ʲ¼_�l�o��e�V։3�X=�
�x��a����A�4���2t��v��n�����o0?h��'e��~����j84��u�� L_s��t�h�ݩ��Ou4ÒN]H�z�b�O�'����/�f'��a ���r?�q�E��n���՗�c)�~�' i