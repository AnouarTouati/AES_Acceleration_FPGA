��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղr�)L��~`��Z��Ӌ*��RW�)!'T�L�	*��s)a���&��!�������d�R]�� ��L�5;�0�~��ҹ7�p�Xg/�Q�9���'N
�͏�웞:?�p�=�Ud38t�9鳬-jb:�m�ʅ�8S�󜣴{�4�N+�UBfH��ms��>+�=�}ٌ���KU+.�� ��d��y�a��,ޛK,��&%E��6�_+�n ��w%ч�i��z�e!L�<�M�fq���-��V��G���Cu�o^��2�A�S��T������e�j�.�k�i+(��deW���'���(�5>0��b7���RL3���{"-��ڂ[Ft�'�5VѰ�|3��a𛭁�Yqy�
�.�"Sx�h*�&������[�f��4l[Ǌ]����P��Y��Z��bXý�`���o�0����GR��'���$R��I���H���8#ټT��@�7�	��]i�K�B+b�:E]�E��o7�C����\�p�>M�ǄQ�p���f_&�X�ޜM��f���I��TÏ4MD�lM�իƿ�Ǚ�w�ӿ�r �6a����X+��T����z:l��s<�>���Փ�%$Х�1Ǿ��{��8����Tǐ-_���FcC;A���)�`Yt}���ϸ�Խ�o�}����L����%`����i5��=�4Ʌ�R8n�,���)��\��)M��F�,>N��۔>�!4��vʝ�kb�pJYTV��DY��W��������'��"� �՘9tC��/�(�/dѪ�ǖ�J�f�<�ޔ�{4���1P�	?��y�s���
��(1o�,�T��\���?{	��G��-[2$��H�M��N���Ծ�/8E�(o�
ߥ���GP�tg��U�K��T��Q3}@"e���2����&��y�LA@2c`����9$��/�&ś�86�D��5���poO�s��t���Č��h��^Q�%=%�jo('����I��C��}�d�s�(Gw��,x@���� Ld�k�y~S�Q6{<Xy�e7١C��k����&&�~���^C�؎`��� ���&��i\{rQ���^ļN!��y�.�d��-tDQt��(d\��53�
��
���PP�K��I���S�FG-����:�� do��Üf}�[�ݎu)��TC��*Y��l4����HĈN��A�!��w���Ղ9@J'H8�p�k�*�@�Iv��xޟ��|�G@W��(Z���㱡4�C�Ό{8�`ŎUW�3:Ĕ��!bB�t�ǈ�i�G�6�Ē��2w ��n���}��D����+�	����=#P�q��r�����Z �}���+��݊�9�$�B���� ��) B�Q���W��3 9���ބ���z�*e���3��
?���5�����$��,OS$9����V7̶�U��7���!k���[l�����{#��F��4��^0Ʈ�,#NV�����8׻��e���8���	߭bXz ^�J`К�0��_+[=��G�T�f8RP\;E%�hM�A���V\uL��tz$.����DH�����eÆn�j��fe�&wq2��D	}~�@rM�X�v���:J��g�������!#-%�Q��v��z�fW���u"�Ho. ��l]���M���N��cb?Z�<���_|��U���G���<Q��뻜d�r���,�
Td�̤�D�Ao͜�u>	k��dR/�CVZH>�R��aI����,�`�e���2V�L��9:�e�8�&�bs1����#���-�;qU��;]����7KY�ˌ�u����3�K/hV�bι#]YӨN�cڃy�7*�Lc�6�o��� �g7�.1@;�kH	���U�%���ɗ�ɱ�6�;쵕<��Ƶ�l��ZX�'��6�IW�Z�ˠ�r��A�GjO޻��[o�i�S�p�y]���m>O�P�y��|L�ї؊Y��0�+�'/bm/���w]��2^B0�Q��Z��'B��!2%̖��"�D۬J�=͵� �FtI���Ѐȓev%4��8��la��1�#�O%mbdm_OZ?�(I/�h���7�b�6�Cp隥k��c���dZ, 
���yp��c��4��U�ӴV*�lֶ���{��������-'k��g�]I������/%7�Ⱥ�Xa˓��CX��q��d����]���X�[��x<۽9;��	����S��[4��7(ѮQw`�f�Mff��o����:�d��U�-��Av$k�}$>�z$�2p�g�7�݊�����ӓ�c�->t}��㉊ߒ�n8x��"d��6B�a����wڌ6�F�Fku��?��v	�Hk��i�(�5B�ݧ-d���!�j:�'��Q+�&��i�\±�Q7� $&Md��8��W�U��=�W��oe]�����n
�ѾL����6v���)k�($�
�PZǬ�G��o��J2�t�`�V��3����I*�ٯ��h�a�
���ρ��;��9R�ZC�u%@�?jL�~�?稀P��7�TN��J&��$v%+!q�	�S[-H�7΂��űY�c)ɂł(#	,dBG�=�.�h������ɰ�-��2�����i}q˚m�&�l��?{�o���D$u�d�'XU�W�����V��pĵsI�<C�N.�����4}�ʛ?���f�_��=(`�� ��R���m�R�W�HR�;�t���Cդ�zG%�S�W7_=P�T;��鵡��9���cU�����w��VVʱ[u^©*x���ȃ��NE����?3&�7��X3�JC�Z�;vr^����Q$�Ve�$�(#j���v_ab�<[��%�����M+�Y/i����9I�$0�6Q�S����l-�[�����\���(�0�s���Jk�K��ƈ,م��5��%)C㦬��ĳ��t�t�m�J6�yfu��� �N�:�;����j8ObL�К�[������.,d?�lصz,LM�|��&QՒ6I� �u�(�8Aw�b�BOo��D�{��@���5�'-�	�Ӌ�j�G_U���k�f��ѷ�x�h���᥁v����4C�|@�8f6�`��s���{52��l�͞��t��
����WI�Ez:X�5�y�'q�A���[~�r���"r�AVv�*����X7A���A��f){�͈�J��?��ޮ� �	�gp���hVw��.�slf��΍�2Z����k�}����^=��+j�ea��7�ߝR���pc�vn���#����ۼb@	p2M�U�@!P���uWN�ߝ��K��`2[����9�t�i��j1���J\�&�M#�d�̣y���áPcX,Y���yD2ԟ㮗���>�2��@���1�����i)��=X0c�%��GE��A�i��߼�P���5�~�H����40�]����"�P��
�ܭ��J�1���狁���!qi�c�9��ee���Tx�t��H���۽<�f����HK�s�N1e =�nN�Gr=T��~<��]ԅ[�oغl	W&W �H,�d�����l
skK'lw��X¢Jd����_]����w���2��%3	y��Øf�f 2F����	��@�G���kYӇ#��ئ����o����;��� ��$A�W�W�\���E��1<pǽ?�ˀ�Jq]�+X ��CIj�6��k�׽P.��`E�y�x�
�ͪj�U�e��{�i�ye��(���J�ĳ���AK�a��	�$�,� 2)-����3���vug�Y[����Eaw�� ���V`(YF�qzQS:�'>*�H-E�,�0�uR1;hD�rh�9�ݹ�J������(iM�+*�?��t�*U(����ZާX�r帬�G��sܢ��4��#�i58�!�f�s�u�f}�¡S��^�pl�F䐶�9�ya�M�T�8��j�j�%- ��at�b������@wh��/�� O�M����H"�\�蕽�Խ(�@���'��� �3��,�@�-ywdN���~{-�����jTo�bXkʏ��+8�wF�wlM[��ع� sy,.�?��P2�n�I�U�t��ߴ��$��5Ĩ'E��*�����0U~�f�L��P�<�s)��D�Oj���2B҂JYnR?�f��B*��.o> {��=l<��@��dbXN� ��J����"��[���q��5�|]( S���%���9^ž�Yϻ�?KB�7��j�Q^ӭܯ�=��`�	v=��� ���� h�!32K?ܸlV�ED�6R����m���}x��忟X�N��#������A���ĕ��uZ��RQ��`β�"��h�&�O!ۑ
+���ut��(Pq�`�GW銇��ϓJH����wB��%.w�.��l�=�6
�_�P�±� �����An%=7HB�@��������F)�瘄�={�Q��ˎڎobz������оl��IBRUL�@� �b��?\��Y����B��p����.�d�+F��hH5>!P��m���^L�[l���N��V���)�o�Vs���GʺI�§D��J���z���G���8b�����#��+�~]A���l�0�Zaء|�P����&$��Q�#��
 Yۃk�����:��?����J���k�W��j;��Z�4�KP�	��m���8�	�`�� ���Ʒ��wBĤ�B|�_1�)An�fm� V����t���4Cw��-PvRiU�U4��yv���0���#�^b>�j��ڿ�,�p�n�.'�}3ֆ$#HPʥ��NѸ�A
n"�����X��S�GƧdJ����l���K�G�,��o쾭�RX�1hG$2;�2��%�O����! S;�3��bd���g�U�_�c�T���=���d���R���m� �a8�{(���ȱw���O���|�7Ů��B�����:"(�ya�tm�t���y�"4�%&���Y^�%� �M�ޫX<�Ƶ_�M�A��{�y�.��|�;��A\+��pGa_��Sq̗���n������c�w0h�ȣ�P�#~�=u��}9������
�g��mLQ����su[}�0z�َ�.������M��[h�sZ�>Y��"D���S_F�?	.Ϊ�mj�,����Z=�K��A�׸�X�'I��RDs�&�$�kSTNcu=+�Bhr��K��ț\�� ��(t����W������<�C�Q��
����q���	�7:,6�-�e�s��#;��x���*�!Ҹ�%fx��n���W�<|+O�	�*�3����E�8���'4W!��Sh\��R8k��'L�0����(�<�F -Wx�(d�8��O�)B�	V��6C�AyV�1P�����"�B?3��������(2$�-��|\|J�˙��Q���3����Y�7��rF�҈
�?W ��f�z�]ő�K^��8����L1���Â�. ��,�w�Y�P��M9"����u-�#A� ���cD�����O�&)W8�&s}�@�0l�.~��X�� vb�߳��<u�	��U)��S�/�_�Y���X��L��㷴�r�l��5�M�Le���G��cKH�k��h6T����F��	_�v�����,�iP��Gf}L߶?T���#������MxO	:Kd�\�U ��A�$3�hO���$����)`�Z�\��Mo_�B:İ�S�*��d l��)0d!Ǻ����B^a6&�g_�\��*�R	�\ ��/*�\��lƯǹi���)q��5��������m�G��ICy~֩0�;`�g'+]�q�r���F��٦�����ͨw;wL娠i�����OA��t�c��b�C���R����ѳ��K?M��#@�8�yG�&+O���5����)�6��%M��C���27�y��G� Q���%�o��~*�W=�m~ϙms�4إ6�d����V9�����&�+����2y^�C���ϲ=ڧ�&�zh*	`�}�+�É��a&�!������fL������:w>7P������i��aJa��G���J��^ƙ,�y&Ǽ�$�T��p�+����/B�����8�ԋ8�cC��Z�[��I��S�h���EO��Oo-[�CީE� Aj��s(���6��J��l�ո��U�K�^E��%v\�>5�d�sl���:�c1�Q�8�4/K�.%(��[�\�2f�Wn�ߍǆ�,4���a)?c�
C9T�
z�^"�e�99���W݂�w1O�&�(���h�$�Z������-�V�����"��E9�>���lX�|�Ƀ�o�l�sD��6���Z|���b�F��:��5�Oߟ�W�H²�����|�:��^4)P�6��jƣ��y��K L�O9Ҟ��^"�C!�*�ךCЎ\k���Һ�n���7=��5���ry���t�b�笳+��~���5�O6T�eaԭsƊ{O4Q-����^��D��/N�}�⳰�V���*�Qz��P��r��X������cb��!*�J_�x���'���f ����*�JR �JD��'���*�m){)>��w8��	L�7���	�Ci�[W�}�o'ܩi!@!�]%Sf�,��k�5���|� ���j̲�[:}�%�g;b\ݳ ��V���_Q�s��E?e!f@̢��(���䁚�Ȳ��~ !�J[_�$�y�O���vG�6T_����]=d�L�@Ot���*�7`��GتC׻�>l˲P������`����rqKj��h��'����֋zP�!L��1��2� 1k��uAwd�����}/v�iӵ�2�4A����A8'�M�l�z���5�7�P���Qb����Bi.,���S�Ȉ�+��γ|f���!��Tߑ��؏��b`b7x�x��u��܏��i<��fׅb�͙�X�
�{DЗ�i�Ю#RLl�O�\�3�e٫��^��R�]�l݅�Vr�TLÕ��1:�z�f�.u'I^���V?ք�N�Y�-��L��WӴ�6�#��4[!P
^&�=�P��h����Ҁpm�J���y��EsɪM4�}�)�ԯ���ue�]1�
;�u��b�6���2�+X<��ݳ�s�~�IQz͓C7�<��0*]
|��<();�]���Ӭ��۰��L;p��Fd:, ���vK��:��9�i��A��dUm��6�8]t�8~�5E[���7Ą�Cw���ED�\fU ���*����4e����u����S�Kx�f���n1A�_��d^Ѩ ����(%�i�7��Q�l��zda�9*�!�W������J�W�/#�x/y�d,��j⻇�-9H�q��/|$�bR�� �}C:#��j,�����;�����~AA�m�[�m(>���cj�Et��A+�L�ݯo�9nD�W����h���Xu�(�א=����a��x`��L���y'�0+b������_����4K(Y�D>����f�q����df^�ߧ�!X4�k, w��K$y��U3:��B�����IpP��[���q	�r��i����R1�z��d�e��*�/�����NV޶[�o[1�m�0����`�L\�Z�����"Q<~�\B��2o�N?d�b�/��Q/�s������5�⋪����.�Na�MH��z�� ��J;}�q�~���{�0��E��z����Hݣ�@�fK�D&t�S�#�tG��8�|� o�;�� ��z}�x��P��&�h�ڰE���6	d�٦W}�pW��Aϙ[�f�ZB����/���xs43���ٸSѽ�I;�^}t�_O:�\���ӵIe���z7&�uĿ�:?�?��|u?t���|'�q����̲0P_���G�c��� h���'����uؾ���/�|��Sk�@¶�E����C~�*� �u}5r,�_�IY8wB�HȦQh��+�۱1�8�l����d�I��&��*o���p�z+"��'���1e{���d�r)��Z8��^���{cPY�l�u|^.H�&�T;~�K��ɀ����XV����~�B��LM��Š���{��p�(�E�/�Jy@�v����Pa�z9�D� $����/7K�z��u����'�=Z�k<J�D~��c�#bc��OP�ik_����y:�����Ԉ�ܰ�}��;���1'�`�=���m;��zx̣(^��y~쵸䂾3-�˫֯R�'N�^�yz�l��4H��~�~����d��>�@�c�w�\�.��eU��?�|�hf���$�&\�q)��?^́�#<o�nA���Z�sa����OA:T����]�����(q�7읣��t�����Lҗ�H@�����G�M/����\ˊ�v��;yXc�%�8�V�yۦ�]C����ޅV/�ාo��GΫ>��?瑼�2���-*BO#�)0}(:)?(\|Ú�RI<���YkA��szR���8�*�
4�Jv�npNn��PR�d{�i�7FIV�hÚ�~��(�b�K�{Ef������1��E��
��Z�>0�ʇ��>�NA.;h���Ȃf��g8߂� '�_�λ\��n�*���f����U�W9J^�*�8�m�*�W���9/-V���u����F�T�(��J��F��KRh�6!���]�0a���=�7���L��S} e[�*ʡ���W;0S�E�ic��$��@¸i b+�IEI�Q����Em�6�$G~�Pp��uH$���t5l���u,����7�[�r����Н�����Dx��vO��%��7�4Q/P�܇��L�U�zUҝ�:��3w���"4�K��n�� ��#1�a���A���
�ad8��b�����"0�DP���m?-I��'M<��eK��Sf��8�	=w����+�Zl�P�z���&��n���o����*��D��5'��jóZ�ĥ�&���Ml��7��r�2Ha���x�����6��KE��0�"�_�r!f�Bv��Ä�I���SB`m���&��� �:"%���׆@��8�����Ug��e���+ �����N��v����p��\���FkG㙳b��U=r�`b(?��d�5Y�RY+��#Y4׽$gHU5Yy&�'�12�4��I�?ȒM�V�(Mo�Pvi�~()���=R��{��̵F8I$M'������O����Թ;=�Hm#�_����e�1��뀉�h3����V��zL1ne���K2��oz���[���_�� ^Γ����)m5�	`H�&�	�`H���c�L̃�Ü�A$$�������F��Ta��Q�9M��z��A�y��[	�����&5�(5+����Ң�l���"$��u��`��?��eE�}�b�H�|יcBة���"ʌ+
ݟ�6S�ʳ>'����ڻk�n�?�À/�Z�Y$gA�W1vq[>Y_A^�T3�س�M���dڏ}�_}+N0�"�������T�h��Y2�{��W�1럏GR���a!��%)#�}{����b�;窡�_H�-������zX\ț���M�N:��k����#7}3�zj��g
%������9��<U�fH�2�L7���~E9D��+I��<���3�r�z�E%�U����W6��ڍ�{�E8�k��_,�ۊ���3� ���U<��<��t��_	�FJ�ݯVzf��b �f��H��=�%dy���c��t�NmB�.+U8�ޘ��G��UФ0	}/�L�1kd�!�%o��{�rCEHG�6Lt���Ͻ@[�{��:S���'����1ͷ�)�����Q�J�e"��	T���cV6to>U7��^'��g�Z���6Q��ϏX�rK��7=^ �_��E����8p��/(�n�,�=��O�Ф�]DD1�y~"}ZO�κ��b�ִ~*pT��@���y�*���#.�u�z	�u�RL �$�9�c<�~��KU�����6#���߅	z��	ч4xS�� ��&߰ʫɲ�X����79W����q���|����A�gG���R_�y����i4�O�H=�d�0pd�o����u.�����ϵḴ��}�<{�҈*;��j�bT�e���}@h�T.{$�0���z�u�	��A�"�����nQ���&��<eJC,�|X�y��9j���icI���w^;�F��1 ��Y�"bH@��Di��sw��a
������I쩆��T��O� ��B��+K�\�$x������d<L˿:@j��� Ԯ`|�\\A��R��!��#>ם��0A��2a��YޱYp�Mڋ�4p���P�F�Ɵ�Ц�؏�ռk�ͿՕ�WW�������b'd$���!����K
�k>D��]������3���؎�?��͍�U=X�%t�^8�!َ��������	�#���:�>�����;�;g���b��eE���������w~/6;*��)׫�ԓ���l+��>��xq8]$��Z�ˈ�I6=���^{c�xD�s��c8�!����+h���E�*�?�z����N�[0ӏ�OA������0 �%>M�8�4�P��c>