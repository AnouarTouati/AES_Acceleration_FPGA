��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&q$�7s-u���RfS�k�ݖNзnU��.j���H�8�Z+�б�"NT�]%���Q�ƙ�ê���d'p������F�*�@�D����OU]�b*D����&�+�J/��%��&8#A��(a{eѡ�N+%�K�r���Bu[������C!�I?�T���o?L��$��=1`��鞍~��|�m�G��2P嘶��X�����x�.��x柉����T�
���M�b-��Ry��EXw���u��۱���2}���D�U�������vN���C�^8M���KTJ�/��Xj�+B�F�T����jY�sFC��X�1������]m�+��i�
S'䏄�B8*������/�ر��z۾�,�_O@,�j�5�<��Q�)�1N��n��)w$�S��5k��lS ��LӇ*��:f�CM� �)U���g�P�.2��`�荌N��V?��s��h��2��<�?�X��?�DnaC�>�0�P� ��/c��~ԔUo�y�O+�k{me�Պ�kaNq\�!v��j�I�A��;�y�O�[�-�ܔ�_3�V�"*h�:Hi�W�l1rL��#\Q&z)Dn����f�i��p��=�#4�����Ky^h�p7�)w�)/�9y�B�v~?���7�d�2�p�V�wpϬe�G�V\;f"r���)���G	�J�r�y�Ց|���(�y)P�P&��n�����.S���Y�����-P��nk"�{GM�� ʵ2�Z���@;~���4W���ht�6�5g����Ճxd6R%z?����7��Ӧ+�;�BX�Iە܈qa����+"{mN<�6/�ؤ[�÷n��Mł+�~S��WbE���mL'��Z�\nY��:CvDg�ؘ	�,��P��t��� �e��[��{����u���9\6r�1������>�֝�i &�蓅�7fgլ��
�����Vx�aE���b46�KRO{�~D5��_s����ީHs�����WE}�د�K���(X��D��hƣ_��8]��+��% �k|��!�$�M���{LE�pZ�'Q�����9~��L���Z�BTJ�*��t���!��C~?��#
`M��"c�4�j��E:Q�6��ع�[�ä��k�M�4:Ԑ�)p���2#j/Vo��HTT�?$ӫc��'��ae�ɎF��2�$*�S�u#�|�F�� +��{'&χt�G�`3�} �'P���+Ʋ�<X��j	��!0a|r������{;�#[�l^;���� � |%�u~S�H��	�5�=n-1㊜��?�.UF���a�� 틽b�O\�sA�㕾��WJk�b��\��ظ�7,_1e����0plb�z=5ȄP��hc�����
.e/�ۖ*�J@С��j�Ͳs���%��oK}�q�-Zn�1)�2^�����	���E5�!�՞`v���\��̎D���h�L�w�~�)�"�ä�|��X�3V�/�~��WK��r[#��1k��v���!%�?{�cdj�i(QL^dNCb����;�����y�c�����J�v�x�S��C�Do�Íۚ�⧋�-�����4��B��g��vy�v��q_����7�n�VX�qY�zf���ή���.MѲQqO>5�_�U6������S����N�a2�`X�]{�S-7��f��*�gG�����w,��gƏ{ފ���o'�>J���SP3��۴��Ub�	p��Ա/�WZi���������68 �i��>��t��Z~������0�"�(��Ά��P�FV�O6VW��.���!�y]Ed_ByE�����0��>D1O ��Cӝ{�]7ɣ�rP�y�D���}�i�Ԧ6ӌ�.S�(�5��e�#΀��J�8v�B�d�i�hot},S[z3)�Š��d.�I���	y!�uV��!��#�%�Y�.h�/�-B��ae�l-_r�����M�X��"m��a,V1Ĵ�0����t�@�c>�J9�&�D��H&�Y�WW�U  ��Y�َ�Şew�WS���)��I�b��L8��gD4-�u%���~`L�p�tz�����,�*��n�� |�i6F����Ty+���}�RN\�i��AY���n��>g��2���Fb�>;��}UhB��G�?g
f��I�~^�y��y����yb۽	�dp5շ�6e܆�vڅip���nL��Ȁ7 ��)�o�)ۏGk�b�V�����V8���k���/ u^��О&�}�a��ն�����Ȃb=hL_��Y�I�������od!PpB������;>��䆀��`=^��#=غ<V���MT1, ���p��ǁܻ�/��Z���̸ۅb��n�}J��O�)$���i�c4][F[ҋ@,�� �Z�V3Î�Mns�������r��t��ەMY���n3AO!){���YA�X�w����i_�����.��]҉�sn=;H�mĶ�|�vG���J����Fx�U,����S7P�J�OD�V��ܿ�ז�F�d�77��G�Ql2�e���Q�X�eơ@z{�p�Ea�� c����u���!{?��E�����el�2�K(�X;2Eុ�/揝f=�j|dY^��ڳ:��u�R���.����2����BX������ ��8�M;M��.�{%C�Xʡ���z��6�~�3�#%�._�3�E���wL�� 3�]k�Y/���f��6�R�K?��`��X��n4V���&���|uXu~��X��׆�)1{�B����yw�j��H��%����x�k!xP�.��O�U������x[���B1:SiQ��{ϑ�U�8��2�vTU�u�����y��u����J����o�� ���?��D["$xҠ��_N�b������oa%�^HIъkʔ`v�+� �s�^T_�Ns�P�-gp�R�c�rC`�Ș�Ԙ۰Y����=XF�"�$�LI�@�}?R^���v]�������n2]Tn���]s��H!b!�L�t����a/�:ز#� #VWʒ� ��J�$��9���K�#m-�#8��e���B����9a�C���ZEM8]eo@�qZN�\e\��p��S��֜����t���}WJ$#u��j�*���D': ���|:��	�7v� ��{�d�m�C7	�9J�[���Mc�]����<�y3.u�j��d���v[?Z�R�q��A =|��h-�jX��^-�ڌ������d���{Bܺ�~���5j�3�N��'i�gl�>�X�bcJ�y .��,��bXNe��(aL#�a��9L=Y{>��*�>����E�y���֨P�c:O�L��o���Xݖ��Q#A��2�	�{ɻ�VG���/���;���^��U1Vo��ò%�/�@E�<�"Ro���Q(�y�?�9��C����5$0��X����3� �Pw�m�m�B�7���5�"(�=�o.!�mL>���h�	?�R%8,l�ϔ�Z�@7�U��y���4q5a
])$��R#՘P�zbpچ4�7OU��0���-��*�yG��{K�~P��v�`Tn�qk�U���ފ�Fpq��R�h�8�K�W��'�<M�e=%,�A`S�-0�J}7詪��G\�3O]X��^I�m�����&���IU��L�+�JMjǕ�G�	��"�8+����w�hB��jw5�h#�GE�t�Y���d��m��Rgx$�F.���[������V���[������³�Q|Z\���+���W��/� {yBw.�6@(�NP���v>��$S�� ��ܣ�^z�ô�1�T���5�SQ4���K]e9!=1u�ZJ�dJȽR=�ظ�~q9����lB7���h�(w3Vc)�)�dQy �0�3r��
M��p��X���w$��Nin01:��ԯ�t{oj���-�5h9�>�; CU�0p���z�x�A"Nfx�ƞ� �nO�ʐFM���@1���ȕ��ng�TB~ �|�-ћ�EP����W��d���ȷw�F,vM�X�����Ы��R �SG@į�)d�l󑨸���ƽ"[$$j���q��e�H�8x�;QZL4�K��dbO�(%}'���q9�L��B1��uJh'��������J��=��JE��\n���N��~�Go�!|T���A}E�bhR��80�ՠ��rP�����׺�ně��2ˡ1�
	P��^����1IYp_�O&nUsJ�;�ȧ���|@�2�P�ȍ�CC��op7+Ti�I��$R�z�I��tH �䨲6������Zg�w,)#N��e�.kx}��W�_���ej�hS�G^q&A~���ɣU�㭏�����uId|��-��n�t�R���[�Y�q���1D]���M�@d[�u�R��(�C{��mH&�NU"aa	LB�>	�k�̀f��s%����b^� ���8<?R���վ��_7G�N:�܇&;�F��Z] ���3�x>�=}�R��CH[y*e�_��0�b�9r���jw��;�l��I�R�͘�]�J�pO�w����s^�2v�ȧ>��usL�W�� *���_�#��V���iBðp�X�F���Ak~~/z�5���[��-�?�%�gc
$�돍���CL[�>h���i��X�k5�޵b���'�ðWY#o� f��Xi����6���F&��&��8�V�&��Rk��. �H�0��w�hg+v-����Q�Gz�%'"e��_=�<���ń�R�R�:�D�N��9��`�>����N���b��]���6���	� �"���/k|9�#^ab�U�	� G�����Ԟq�O�|o�Z��j�J_��.R��I�<f�?�ՠ0n����-�0��P5�Q�����G�����>-������h��j���9��NQ��^��q�o��gϾgw�U}MwJ��*�v7��5-~�]Va��U�"gv�}n����
��;	$JVD�u��Y�����ӳhA����=�[5.Pl&er��(���~z+m���,3������gU'L�إL� r�}^�b�
������MNaZ�U+Ů�N���OQ.�8�S �ʈ�>�\b�&N��y��m����\�B����A��0��ec�o ��ه��T�v<�skµ�Ƞ���Y����:5�<�����L�H��3X���IC�w�I�!����e���t�^Z�1��U5P�e@��⸗I� ����T(�p����W�a
%XSщɺ�3Ѐ��Ϣ��<��r�P�ɡ_a%��_,��b��D /쬵�o�6{D:m�w�Ԩ��l|�:1.�B�2[�G�iN�f��Wat������5W�����_O�_��*|*��Og
a�C��z���x�A6On��K������ι&����%��� h�I��;�_�p��.�-�,�򊗔
�u���
Z��?�䮣w�/�_]���	aE���h2���Լ5��؁'�G�AG^��~���������ݜ���)���\��n�4 �ɢ��
*ji%�wb2Ftź%������6����ԏ�e�_��pm�y��D�>z�U6w��~JUɌT��uA�Jl,�{܅[��!���=U�3�Lƀ�V���)���������C@���i�V��4�;)��Y.f���p0�5�R#�*:�v�~�8I�����m�7��^����V�"S5�Ew�H4ח���}'�J�ğ��z�0S�����o����N�������
�|�s{���IyZ:��i[���U�3�Z����2��2k9�A;����RT����~�l�|���3�k ��������n�����^��tI�IN~�f��2��%��������}�/�q�*Q��x�).D9cn�hu;xNz��O���2½�	S�GH��>��R��G�cS�oa#��Ǫf������!��&Cql��r��	���̌����P)L��B�!�O��X��(3RI�k&��U�D�=�24�޹
CL#�2KX��Tp�S'm�G��e�MaL�V��	�N�k�=��P~i!���^�qط)��1��ó����׵�\��@�#uT���:5h�-vu'$�hB�i�
��f��?�<�k�S�x*����=�}2kT��0����Cr=t,�f��/���b�4�;Z�A�������{�3ƑN�R���H"�g}z�t�����)v��l��I;r��W�m.�JT �j��bx"��-C4E�}SZ-:{JA�:�=�%�#8@�B�~����r����r�����HOCµt�!�Y�T��C���}^�T^@;��oQ�9���D?.�8�V�xq���~�l�f���"��E�nqo�LC�N�����]1wR����6�{�/t��/£�n�����W�R�`	��LL_'̷|��B��9-�Z�)lŦ��v2vz
�����mZd17)!�H��s���}d擎'���X���P)ͦ�"S�о~\�M /�2Xݔ=T��D����f�`�6�`�r �8t��Y`��C�]�_��2���G�3���I�Jo��=�l�Ʋ����tRY֍",�QM���1��/��j��T�}������fkQ������H����j:�|�n���"�M�zD_�YmQ�)�s�]l�m�"a��JՇKca�{}us�?W�xi�k��'��ȡn�Ƕ튩�0�C0�����9�e@M��W�/�]�Z���d��!���]�^����@�vC"0�K��Y�1�lѹ[Hd���*������}"Jٍ9П��a�$iV͛V�,�b�G[���$��u�|���3M:o�]��|�-z���<OV.j�k��y��jJ�l\���EO̚Z^ڴ��W�t��B�����[<���.W�R��?�	;�:nT��0ԈR�7��
B#�v�,	�	��;��e^i�1ec)O�tk�&zj�ڰ��NZ7���3����n�8�<�>� B��T&����)�qA�����nS�P[,R�K�x�։�ېm�[�#�d�3�_N�}�l;Κ�/����Va�7*���լ�Z�I*٣_靅���I���+ظ2U7SoR��f0u8q��x�sc�`)�t{B�51��3
�%�^��m�
9�ͯy�'!��^�aPѦ�+&�������k�J�}~�����k��>�S]_�e�Y�@���e0lA}���&���i[L޶qgmY�v�U6�g������k׳�u��0�1Ps�%��p]Nn�ҀyX��%(��kjp�饃^�l�A�%��:_�Y�9�[���5�;��k�&��h	FU�x����w��+��
f*n[����9y
Vq@��$��|7�L�����	�&��kaZ�sI-�u%��c�:YR�pƄ�E�!5�ZA# xc�4��
_0R�MZ	k�ƞ�����ާ��5掤�n"�aY����x�{�},�6n1�'*��&]f��(��$N���!���r���lJc�oEK��#�b|QH��v(�$�u����%}���<�*$�i��tj�.�e��P��M�w�˫�Xҥ��&���֛SC���M�f�N��K�f�J	�Z�	Zsӧeױ��^���'_F!66w�k��
�J3�q��~�g3)ٰ�m.D�2����zA�r�vbz�Q��u;B�c"�?��E͟,�e�E��U�Gr$Ayk�G�ֲw�TK��Q��HP.����ډ.�nO>.�����ҝ]���=Q�)���r��U���;�<��4(h��7Ѧ+(�O��f�}��\��i�`]��5OI�2�ޙ���"��r�}��1k�� ���>[]C�h;���� ,��$��bc�����C� �- ��Ka4g�Cl�E�f��C/�l�>tU�o��2ν�g�����Y�1:�Y���z�ha�7����$��41sḸX���5��E�v������[k��49���c"0���jV�0�2��-}�)�<��l��܉����{�y�����̒p%�Iw-9틁��p>q������dՇ�`mS~/���˻"F�l{lgg���OoΙ����^a�|,*g�pEc(�MpO��=Gs���D��^y�O1qF��j��V�\>i�a4U�u_%c!�{�,}�1/������e����ȹ�#�f��3�h�rTTS��	q���;��,@��942HI�A:�!��q�V��.���E݃Tn�tU�`�Q�w\���auHac���V	A��E��V������$�.!A�S��e�����H��^@)"���oRy��ι$��ॺ�vN�uU�폻��?���Hm��Z�=T�5pqn���p��dI��)�΅���!K�j4�$��"D,�-{����vM[X���5�?v%jc\��O*��	Rҙ/=�<ݔ��D����۴|���h%�c�<�3`�����D�b�m*S�ʂr�1#y��Vٙ�G���@P�8�p��xY��m� iuwH(`�0�=�3xi��6Qctv{�&�ḅ���-���Z������,�-6,�Ŕ��T}e���o,�c��㞸R;�Z��!5$Q\���v�5D�U�(Y�ϴ�e�	+�=��a��7b�	͔i�տ;�싃�q��d��Y\^�)q�Bl����I�8��qk}ArrG�s�IL%O(+���Ԡ��'���h 
�TX}��_��Hʚ}��3���	Zc����0�G��\�.�Q,�'W�}Ӱ��	�p�Q��0�nY��'�9@_2$ze�U�ᾣ��U�r��L�"�'g���%��[�smY�O�/%��sյ�!_��&�2����++s�"��}0q��y��:�[ȼR��9�Bd��.W)��� R��qӍ��;ynAupx�<fY��7ק0�א��m'V��O)�����H��} �$�`���j�9^��5��`���=�iZ��y��&��q#����s�fF�Iy$��;Y�WH:�柲,�ٓ{�Zڢ�JD�v�QH�2+�<N��#�V����'��e��l��l��d�.7Z��1��Jx��e__� �Ȼ,Ĝ�J��m�&5@��;�	U�F�B��O�7�?B��KUoĠ�N�/�:������&�5�u~ެX�B�t�[J�go��2�SL�f�����^��Qay7�,7���@��L�H��jǛ���������;����6F@;+��-<}��܃�t��W�{��,�����3�]D'�X�?/;�.�k3gOG��o�7��!C�o�GU<��EF^�9�Kw6gɜ��|����#!T�p�w��*��--�EMp�Y������"ϽG�\o��&�;r�d����)C�д���;�_邲����O�Л�- Á7K�����I�C�<b�׸z��P��AB�Q���9
y�!��߆���J
��9�>)�+�Wn��A���-��ʒ������=�kQ�[��x���);��8�̔D��m)����}�bC��,�9M̟Ї ����MŶ;ݩ�=���j$�1���ʖ��0�1#1H�д5&��('��o,@�y� γ��r��smo����H��6�����̇����dl�0���R�Ku����/}hrF�f�xM��#`�K&�dMqU��4��,�gt	#Tܒj�P鍡���c#p�d(\�
�xo�?F+��a����a&�n�w�,	��୑�?R���=�3�0�G=�9�3�R����Q�Lr�͹�V�+	�m�M�]r�.�������/�.	���n����_[�9��ɤ�5q�߼{�����O�j�sP���`� T���%Ɩt���ȸ�f�1��p%��&�d{�ws,p$D.�	�UD�dS����h[7�C��������͜=$����;�s�� ;�ϫ�=��u���K���IkDݣaN��Rf޴���J"4*��q��P����&Ncn5K��_j��ǥ��u�>~C(���3]���T��.2
#��l�v
!Vޑ	t+�J�-��<zT:����v3�b����كZ�΁64��H` Щ3�,��2^���b��O���ֲI�&ա@ l�(�HpҺ��;���_*z1�\�����&�M�Ǽ�!C>t,AT�O�֤��Kc��_^���o�0C�=���Șƣ:a�4�Z�����˨�lI�pf�B�Y�d?7i�s��מ]cĮ��K�?�j�y�����2���e�� ���'���2�7��S��M1!�7�O/v-@H��4���dN n��7��I.�
��-P�"F�J��H��P���7�R���k"�К�����6��l��G@�l�1_�V)������8sO��E�C��5M[6xN����l��'Y4Nwq��'�;5��*��K�s��:4?X8���%�@�ZE�vъ��=��:��.4q��r�f'3��Iṃ�<��c��`����[�qY�:�C�e�|��ĥ��L>{�]��������'I�⺍�)�XF�Â��%(��B4:áƥ��M�4�� m��Cq:���O{B�������K�tF��o�%MO���XoM�ܓ�-*����tR	��!:�A�RmR�,�r��Ƽz �����ǂ$�~!
���'�A�-��𼦶��s� �KU�����(,�X
8J��81��	��1�4s2��w����N2�kt�j��xt���p���7���ӫ�!%�oD�+��c�>� ��p$Y��l%˙��}�)E�C�+���ъR �==���˦�}�2\��7� �\euAZ��ɺ������/�;�p�A�Ȣ���>7��YnU9\X<'�nz�d<�i���%A'kh��g�qaz������L�b3ا(zj��9����zQ�WD ���i�Y)t#�`B[������ʅC���	o��[f��d�v��C��S��i�$� �I��R��F��V��HJOӈ���ʟ$/��X�b9����u���1�+�헤������4�%�NDԏ4a�2��[m;�=?ze���p�;��B�?ު�g������+L����Y*��]��"%���.�=7"��gŒ2���ZN=�?���7P�6�Y1���>��2`gÍ����P����6�"��:��o��s�~��U"M�1��G�q�j��Nsp���L5%��,�rjg ���S����r�w��{��t��^gVcܓ�!��*��\�$�R���2�K�`UI�����"U��=X9�$O�`_�´Bj�1�f�$uy��"ʇ6GG���O�n��ϒl�i��	wu_������'q&B�?w�bF�CU�&�Ӡ4)�G�h]�����}��F�v�sD�4d:�lG��7�n�oNG5�� R�����>e��!t�����K�gC{���R7�at`���Q�����	rW�3J�3ۀ�)�|�%�Z����>�kPיfw�/~���<��Șf&��[���u a���z!���9I��ȟ p�bj�L���t���vv��5�T�5�>�<ޒ�����s���
m�v��2A��%��kD^ϰʁ���]��_�X�ĭ�0����O^�Bӓ�g5y"��aF�f�}8C�sPU˗4h�@�s�j*:<ҙ��O5��
`��`�cH� ㎫$jr�B�). ����WǢ� �@x��I����Jo�݋����S����� i��rm}�@>\�a��|s��@S�<�M�2�i��. �St�+�a@��6R`�򎺦�v���j+۹7����os�u�g�{<ֳ��ON�E�n�&�Ѵթ)˄�mouF1%���7GVB��ߑf' �׊Y�z[��fӲ���h�^ض�3��1>�Z�ۑL��cg����D���8�h�cūs9\�����v��Gm���1bWﳓm�^k^吏\n1���O�xUUwӐ)����F�WǑ����U��q��߻�_�X¥�\�s��,�)v��K�Nd�����KY,c��z0�P`�	�8L�8����!��cgO�����<�&^�S��ci�;
��;r�����^�qsI��������̐#�u�m����a:f��QԷџ�fO,�!`�^a�,Åe���`G'R1�����!d�,�n��إ|3ϵ!���4r(v�\!�Jm,�^�����X�T��Y��5y�kS ��dG���Y7���cS�L��؋kj���Ųd�	|H���g�o��K�)IN���>^)*r��U�.>��_��G����s/��_�s2��� h�C����]�q�����i��Nm�g���[�rW�Ο�����6<G��{Po	(� ��	ؓ5)Y�`4%؛'q(k"}<E�#!�:,����-d��e./4��31W������nD!���7/I��or�4���B������h�Lr��}������QRSD�F�9hE�>>��� ����]c����r6(�ݷ����dsuNc�V�G���[W�l{D%�'4�r���ak>�~T��bP8�����h)Ǣ+���v����y���[�ʴ����P ���y}sF�zۋ��2֝�aA�ݯ�y�mã�lU�~�+�^qN�UTm3U7��T��\Rs�Di��8�Ř��'�@Kgk'@+��D��HPg�!\�� 6�X�^