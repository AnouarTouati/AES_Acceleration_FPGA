��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P��/�͢��u>��b�]���K�_�cx���A��"�Q��pMl�jh!�G�߄y��lv�@;JnF����HG;ݤ3����NL��[|$[�U�=�}�ċ����;�BO��hy��Q��=�i2tC�r+����"��[�`n�j��A�gb���~��3��lqF	c��y�z����|�E�`���d��ϭ� �R�b�L �-����!Q,ۤn�i���ۤ�Q�Dqo+��sIe��fӦ������8RR�q�����S'�eu���c0�%㱤�:�R�T!����n�˾���=���k�5�����ؑ��gn��xcy	�[��׫_����J��7w���E�W?]h0їlpx�)�R��G오^n�w�:7]�M)�p���|E��#:d��_���e?�20]{��o
k+g��q�=⾰�%�ٹI���xyX������zY���������8�����i$�}Ovr5��!�_�ʣ�>�;
�(�K{E�QB5ؠ7	 c�Ύ���)�Vw~r��|e$]Д�E��G���1�q-�W�����8X8ԧo�;��LX�3���e3 ��,����l���/�sp0�ݺU���1+�fi���j�������%(ν ���:2?�!1Ll���� ��e7��Aa��?�C��B�nl�E�"s3�G��5ח���+��$�L2В*h�锊�/�������3��Q俢"9��[�H:V>�N�	U�[�N*�$RhO���I��l�j�IR�8���uI-�Q��۷,����΄-�S� �t��u/f�ⴽ��shJ��؟�B���ś�'�Ѝo��& %x8��[�4 i��n34�)������	_�� O�nB��O�\�_=�b�oW�����U5B�c���A#  $�+p" Hc�a0��$����S/i�C�s��=�������d�5P난��n��s�D���:����"�qeupb4p� ,�o��KU���sC��W��t��ۙ>n�mޤ�ĭt3r���<���ɨh������gi;ۚ���I�-|32���X��LgΣN�1j0�[V!��W��XJ�dD��IOG,�X�DgFw�y+�7���އ�ƚ
*�SC�Ue���I�"j�rN�	���s�z�X�/Ia.��~�KK��Ȕ*Q��㬘���o.%)�>S벣#Xt`cS�<�U�CX�����L�FBAw�#%�[��ʰ��\��Pɹ��Mʳ������,u��� ��)�Ҡ��2�b/�"�{�;��#��l�3�忀d(���#Iƴ(_���b��6��,���8��,yr<Z��z憍1��K�n��q�L�$�PQTh�����'YOx�2�r9{�qU�����G1v�Q^j5�8�wy�!f��KE���&Y(��/�i7U�a�vF�9���(t���X@S��T|���G/���<�(�����i����P�5��zu������ދ�6�)_�G@[:�M=�T-`'Z���R�O@:*���w�����������.�����mƕ�FT<b��r�K%��!�B �>jM�]`�(V�M�.������F�ȍA��l�TZ��+�Ժ�O�j�(�=�vhG�s<spu\_*D��>�vg橜��r����v���F��7�JPj*��?���/��/��hL+&�_N�V�BL�h]�X��$�p��TxهJTAђs�>Wܣ�H�ʺ���]��I�0�t\ F��ѳ��N��H9L�sV5�9&�4�ȩ�[���#YQ�����X[�5 �IΙ��0�c����l:�Ϊ/2�g_��5Pl�؛W��m%`��n�~�2,�͙{K�l`�)�8�S�:!�N��#�W��D&I5iҗ��F�����4�^{�$��g��V���[��`�3�Y3�Fb֪ځ�*[��:U�c݆t`
����n�|5Dߖ��Ez�V`�Pv�%�����&�K7��gIl�ڪ�K��3���vj#�C�l����'a�~����Wu�x3�!������ӛ����Ŏ�z�,l�CZP)�3��JB�U{���1;�j~��-;�?7�5)�����v�L�m���f��53� ��R�tfXB�K���C��ļ5��u-�I:OmmAr�,�� -:�zr�Yɑ�dj�pA����X�����v�!��P�5�	1�:�eG��S|�^�qz���v�(6YX{��:��A���W��"�ነ�2֗����&��"v~^��kZg�AڙZ���ע(Au�!jN$���kC�K����@�P�ڒl\���o	��f�0n��f?״�K�5u�[�AB�	J�%��2a�Q�#DDt_xA���\������=�9�ȏ3��T�~zRG5U�f����2*��g��]��
��������j[���'m��������U��Cwtw�fz��(�T1�F�V���f����3?�@6��Mr�h+P�uu��^)���$����e�nIE4�=|�tv�\�L�lч�m��c�w����\6M~���}��@�0;�7�w�ڷ��@Q�lӮ=r�Kf��[8���c!�H���}�<�$E�35ZI1�
&4i�$ӄ�Wv���b�9p �y

j��s�^�NA
���ʹ[�,�r�0FE��d��N���Y߿GB��>_�$sR08f�Y�a9㤳�y�z)Y��Q�M������'���=϶k�ug�h�Ln�o�Zɮ����Eh�č��6+�Fd�n�#3hr�i1�>��e�6\�`�� �{��8���뺀]~�B)����&FL0���7bw��~6�kv�	S`���Px�6�Y@!�Ă��H(mH�a0��"�b���j�̈́���)�����,�ͥv��:7!��F
/N�W�=�Zg��	�I�be�Vr��������L��3������{"5�v�����-}4qn�W�Q��1�s��QxWԟ(�;#��׌Wq�D�p%�U�hVd��A]l/���(8�u�6r�����#g9:������\圶k����NR.%��)Q��U�\�p��F���R�J����P�@�8����
��9k#L��}w1����M��5���p�2nY;��L���]�6w���O�7�Wt��lN�d��e��ǣ؈|5�0����L8�AbI2_�M��܌�:��Zod#>)E�P��&��*i�7�tV�k-�_%m1�t�b�d9�	���G��`M�1�V�������z|E�ґ��:� ���e�&D�v �۶���c��چ��S���1:�
�2�}0���h��$���{ nF'Z�W�gp�D6W]���O�ƍ��~Z.?�Si���2-{n��S�+ڷ�X�N>��,2D2�)}������(�*�B��*䲣��~���� �#2�}�o2=����!��^M_��RR�k0��&p����K��ڈ�?�/���a8����Ф
;;�i�m��47�TP����x����=H�'ԝ���xj�꿑����}VHjIeO&M=�V�`K��n�)i�dp�/I�~W}#�I��?UQ؟��
ZW�.�]o���m|4
�oPE�l���+�"�ތ���z��zn���x�'�^��ܩoK�I�-�:��N�1�CF;�W���}��O�.���}���1u� ��0��9&���E��y�1�+��m1�N�#93�/Ƀ����r�w�E��[�y�b����J�F7{�
"-�������}Y�l$2��a��!=I !������_�ן���{!o�~."�$�t��2si��E���ex�(���p���X��-���6���[.���~��d�3'O�]�(��m���x�� ���1��0 }Y������6�L�z�F��r��{?oկ��'��>kn��@�7�X��Ϭ}�,ί����m����ń�A��B+X��`�]�Z��ƶ��仂b=����g[1�aEB��q\T ����+D�Gc2Aiq��<Bш !$jb#��K�wCKK��]�'��00��5�ßZU�B/P7L�3	���4���fqz�U_��Y������Ə��`�ܪޭ���`?�6��
|�N��P%�ce|��_T&Ath4��b��Y�xd�
�E^�;c'�N/}�;z�Y�n}�0�U�ھ�=�9p�rZ��S�I��Rm��"�P&�oPV9�HϬ����9�����g_�:��[�R�'�4���+4�x(��uf���&���c9�kz��M,u���n�3�N��	��%�ڛ��˩�����BV fgm�p��;T������	��%�3��R�`��'��^�r��ΩYcB��_Γ���xu�U���k�� N��|k�����0%��`���0K�,�EZ�!^1�wû��"�}�Ϋb���a����=xL�w��B���c���ѲGB�#:�߽O���oI�X�\�@�Ŧ���I��tl0�}Y�Bc��`d��|�Z�e��Rf��m0�-O�J���#��X��C���\��u�ieBr��@gu���d��[�RO�i�s?��k�Pj��Vj�1�p&��0�jֹ��r	�d4sxO����H#i�j�{�N�7!yw��/�)05��1$���=��I{fd7
(6��r��X��F��JC�2/�2�����}<�+���E���J�)���1R�D�K��u�k_��#�� ���{���9�*�.�v1I3�M�9Y޲��Sk";^�J��s÷�$(w�qB�pi�k"�����l���'*CT��;�Ȯ� ��T���h��1I��lq0J��*ʔ��X2XE�5�B3�Oe�����B+ !1�Sa��H�:$�T�#\��{���:�;M�q�ݦ�{�`��5z�wp$�̮x���ڹ�m3:�)0��H��;*�'
I�B	�ڰ&��yx����nZb���i�^|�ċ��w��qW��r�P�x�O��|�K���YK��x�	39�u�1!�s�?���G�V�Wn+��]Y��� �����>��4+]�r�r �Au��Дy2jP�=D��4lh�X�Rx�D��Y3�@��3WjV�?؀%O�Ɛ�P#H�ΞV�r0�js#1~�f�T���'/AEFݱq�e���)zC��]9��G�+}F����S6H\@Y/	�X�q�Y�u�*F8��.3 r�p��+����c�c#3l|Trl,�����#�Fg>u���\��=J$�o�˴�57��-Z����D>sUt-��sa<�	T��XoM�b�%��D���;�S�f�!� 01�NǐXq4�CIEk�l��7?�<�K�ATv��%ؿ�d�C��Ś��,�._t� ���P��0$|�ur��RɁ�Z�A��$�� ��Fd�@�o������]p���?Dύ������cGB]6���g�'��nS�  �5���2ri)cn�(q��~Z�I7�>~��9u��E~W�q����:Od5t�f��s��{���1)?m��):��2���׬���gq����G���X���{ٞ@��#EYg5M�+	A�L�=R1��仕���i��] ���#�R��a��{���I~��v*ˣ�*��?� k�d<a�K��
3�L�-L���v����pe v_h:q@Aj�7$��������	h���)��Z/�nH?���#} `�7�tߑ�9f�`i�U'984�i�,F�XI�u��pVB�jě�ڻ�,ZN,�pf3CI�k�G^�8���:m�حώL�i��sSqzdmZ�7f� �pD��W걭��x�5&YiV��Zn���*Að^��.ʜ�Zɒ��ߩp��֓���`;��ő?��ȟi\�Noq����o3��� �|����W8���|���ߜ_��1�F1W��6/��q�Ӡ�1���ڶR�#b7(���.��"��2Eu�6r"�So}�9������<�[�Mz�Z�Bf�Òf�UI�t���'UӅ��*�I���q���	�É��z�?�0��|1�I��(͢�E-~I�'|�!�v��+s��.`ٹH�����#	,����R!T~��3i�\p��!���AFqd+�?L�x|mΰ��T�ۯ�!�_ԇY��%\Mu8��}61*q�[��UKσ���	�hp�����k'[��r�piP{W ��Oүg,v%a���zYx�m^��>@^;h��~iVQ�C��Cr� ��Ԉe�32c�;�G\n�ڗ(u̱�Nt���lk��/*��^z�,y�e��զU�N.�r� +�U��Y�1��x�JZfP�b�)�]��\���j�L\�"t+ ���#O4�HH7��T*H�d��}E\TG��=L�ť�[�э�Z�
T�\�Z��+��!�ޜa#C��Z�x�B�e���㔘��_�'�%��KC�]^�%4��Z��$uP�6�.?"J�H0�Q���/�F��U9*��14�W&�vnP�=K��jfq��l���_o��<B���a�Wzr���rEQf0��K���!7� xĹ�pzTC"؝�cU�$zR�UKR��KjG(&.�@\�.��*���a�5�\!��?��b���v�[�XRݬBY(���*�l���KD/5��X@܋�^ijs�7�k�|Y���Q�|B�?6k�����7�HƋb��G@�W��Xj��[T��s�b}�bF� .\q=�gw1D��ڸI6�9",ܫP'����y2�3x���a[oC�����3�=z���x4C��*Ԏ�-]��ҙST�@F��r~ß��`�*��J�!s��o�"u�(���Ax�)p��HN���Cio��9����~�H����t+G���T��ϻ���w�nY[+��o{Z^����c��^�( L���v��ݯ��x76��}�>�U᭮�FD����b�3��i0��£���I'ݲ0�ƕ,P6�)�@MuO��фo�
�pƁ�gI�H�m�^����m&��F1i��ɻ���b�J���D��n!'~_��x,?� �}�ZhE�5�=�1�_5�$��`3�_��^IX����Ȧ��ƭ�u}��t���}��$��O�K0|�ո��1˔���}�W��88���PW��|��Vo?�w��t8�a^U2�'���1Ю��(O��r�sn6o�|�2D">u�Zz��g%晧��Xꠎ�c����J9a�W�n�b�P����aLu������{�4���XH���	(4$dr����{�z��������/�l;\��Qw����_utp` �v��I�0����i�M����lU]�zP$���B�`�]9��/���[�!�G�pC�"�,TƎM�&��Uؓ1�������){����a\�cЂ�3�$�^����u�m�9�n�	L��a�9}��A�"�v_�@�c��:�هZ`��3a��kW%����L��#W�0�|��&�w_�����.C�;��C�/Ŀ�$�L~/$ƮWd2P���P{��֢o��S-���s�kG`Gv�s?�]�p�u����H1��i�M��'����w����!3���.�,��%�?�>�Xb���A�ӱFQ����6�I�u�Y�_�
	�Z���j��{�D�{h�&
Vd*B����f\��P8���e]�5��JBs�T���HW��;6n־������	�����k��{�Ky�A�4[�/�"�_����',\���:4�/�[Ljb�>������f-j%w��G20�EmQ_�ۘ��y��S\}1��w5�= ��
K���!�����])�6����J����1��q��4�rl�P.�ʪ��4�k��D4�kuٮs_G��w[�5[Ζ��#\
%�//��![Y%O,
Q����n]�I���Q�([�}.m2N�M���!����ِt� ���&+���9��S�:�F_7n�(��_�7�Ga>���_˧�y��$��KeH���!v���aە��$�@�5���/��|θ\Q���n�yF�;�By��)���vr%j��֢Po��y����c�#'��r��1ȺJP,o�Ow��.�I_���8h;�y�[4]���L	`k��<��D�>��Az�� �[jŪ�r[��5��8�a9ā��b�,�Y�����ʞ���D���������!S�xh�K��q�0Z!O	��R�uH-�\�{�U��0+AV��m���[z����';�4�Wsya��ql�����цBeb
�~͐�̵@E^�������B�w�q͠��V�q�cq�Ⱥ�Ah�(n'B��cG���j��Q���E\�*��yK;[
�n�(rA��)t�)�N�&_i�kA]�U��,�iX��^ ���)~]�	?].�%i>�_�[��#�w)buP_�+�wg�B�0�;�		3Z��YI5��`_H�|S<��H��M
QJ5r�:���3�,'~sf�1��?x����u���YӳkuGX/U��������xFYU:|���ڐX��3�&��ZX���H���c�����m/%;�<�_�c&��̦� �!�K����.�쁺$<L���y�t}��Ao׈zV]9��d�b�}�:��J<�/�5G�6*�e/ �7C���2>����=}%�[���<���!f�_&_��c'��q`Fr8�y��b-�/Wt���k��#�F�TpN5�B2B���0įĦE�8�ֶ8e�fB�b]�Ǎb���4:鰜 �:|9���m��Ƴ~�q`0�CzN�V�0�	\�#7�`/t�z`ʋ�L���IX�ɺ��>�.�]������ܣ���-�a�&b-�R�,ٯ!���{h�6��P���S�g��jm9������0C�S����X��V�8��������ϛ�T��n��ML���w\�Q�>�Tɗ3�����_rH��R%�vi2H�Ebi��BJ���������e� ����%�B�Nr!;����W������J�^�]�o��R��qP�&0�I�)6p,f�5<o�n���t�d�}��(=>߈��J7�C,֍Wqa��1���r��s�J@ �A��w�@i�7ϰ�=�Q{(}~�\M�[���	%B��ֲ8z��c�q���/9D9���h�r���疣,���1֤`c�@8?Q�GK��Z;�-SϜ_y��m�ּ�W�p�y�?Y���ۇ�Oђ���^
��&�Y���/{��e&��0��dk%�$:&�+Έ W�n��1�of/swJ����8T���5��+����e@|!��<��+�z��X���xiO��Ԟ�f�� ��*�Qm*�/�*�
t�w�f�Ze8#Ņ����c��AvfD��48��H�z�Ǌ�:`l*Qv��>WkPK?�B�N�=��~{�欣���5t]mNO�����#&6h!����	g:���+��e܏�D	���Ts�Ȏ�0+-B����:2��l���4s۽�Xߝ<ȣ�a͂�񊙙�a������YBd>ah$�6̽8�� �5Cu)��hE��z�n�pT��)f9�zZ|�
���֒�����#n�����C��^�IO3O� ,1���CdI.���������h	a��NXh�b,�J|:!l=�x[^bQCFs$⟰���<���ĕ�!�lWK���ކ)H���v2��սn�o#7�q}��Ĵ�ĸ����k�'U�mQ���_��y~�U�Q����~d����E_$��*�#����)�X��ӴJ�:�`L�&��Oc���?�ڪ�C�"���vw�|E4��!�U��,�b]I$R8�X΁�_s��Z�c�y3�R�X�	�!� �>T� x�sԖ��K⮶#���Ll���*9O-�!��n}��A���b=���9�� ls`�)�8�K�
�W3��@,�.8|�u� �c��?�0I3���4���g�˝�q�s�P}3v�`��Q��(z�ߚZ�1ϝa���6k�\l�o��r��z����P7{p�ܛe���M�!,ȞoV"����| �34:��\H��Bx��%oIvWy8��9iԼT��o.�b�T�)�m���b�A�@��A�?��-'[��C47g���	d"��*n��G�a7���){uP���ס�ge4f���o���[�n��/������`W��F�Y;&�o%�q%�U��v,_�CE��~co�ň�y�����<'����G7��zԬ	����b���5�r���T|Wem>��N�K��6#O��C�A2bk-�ӝ-������FޢWWOg�!)�hAZnrH{����tG�8����=�9�}����.�]�+��n��O+�#u-���љ�9\c�����cw~8o5�f�?��֛������(�Ï�	�V���4"c=N7�R�D��� �ۦ8c8�)���E�CY�x'l{��x������l��֊�Y��@�~���� c�ؙ�g��^Yɠ�?�c3�!!����P�+�(�/	3Ԩ������@H�<o��\��TR�h5�*t��;͎M&cBDT�(-��Wd��!�
�<� ��t��S�+YC��4�ӫ:�	=j�|�['��O%���'�OO�>.3*��� �ںat�nϲ��{��Q3D��m���^���>G�����*_���ѧ��Wi�]GJ-�_�.I�{MJ�-�p�_j��7��'ezy��-�Y��Ԋ�Cn�LGw"��$�
�����	�fdX��9�R�
%�uU�d
X�4 �98֕����xd�	r�c?�IL,�������
�2��Fv
�V\�li38,��;c�_�ĐG�naU+d����������`��˕lPu(�o��@���>h�?-qcO��T0�^�C�C3G�ݼ�҆����(���'Q>k�]>�;����Wl2�67��X܈�ܛ�e�����(���p�ESB��F��TWO2����S]kl���$�f����I�3��U�1J�H�}�l������O��p�'.5�y��!��y9�L<Ǡ��$ռ�y`�Ĳr�Z�I�����I��y'�{�+��O:8�P5��7��)I����CmT��6v��EO@������`�rx�yC�:xSc*����v�0�;�q��\:��� ��k��VSn
�D죺B�m�����ge�mǴ%��^1Eԩ�ت�v� �	��S�ba h��8pl�����Dhhme"�Q?�<��[��R<�fɮ��ل�|�r���\��V@�U�S�?��1��ъ����݆Z�_w��ـ�O�� �w��`8�� �&:H�4��5����7�ƚ��C���1����l�c��j��~ֳC@s��f},�U��W�o^J/e��u�`\^�X��c�Dn�	�T@F�H��3T��	LR��(tRa0�&��������� ��~y���p<�Aj.5gN�'O����L�{�LI���+�N!2��j4;��/�_�woH�g�һ�*�%�Ӈ=�נ{��7'��s���?��\C�`t�2+�J �
���P����y��ìq��F�=2�GH������z��`ݼ1G�G��u/�u��]�ﰕ:�Y4�.=4 ��*TJ"k��1U�쯘`|m�:����S�^��{#�VӸ ��YB�c�� �� �M�ahc㙳q���C�� �����LA����dֹ��o'�y�������J�b�0���	[���g�{��#�]�`��i9�l�ʥ�ڞ��9���b�aO�cU��K(Gq~m���.�Y��6ﾈx����5n����q��NE��,����9�.������Y�YH�d6D��a�f���FU�y�N�;���&��5�黢���5u�v��Pl��Y�� �E��A�1M��z*��0o*2�>���nP0��WA6!㇩����ۮ�����m��b?�WxČ��XJo�#�R~ZwF`�Â�k�c"�ڇ�?�my�ϋxn��C#��]�f�w�O�F�������nW�7UH�E�	q;��r�o����f�f��_wA��Ju��tO�Yl%^L
Z݁1�3�=o@��2"7I���M�n紦SX���&�(<A���t,�誚���='i,�8��g��?��gc��{�ѻ�5����ZY�˨X�+6t�	V�'Ȳw��d��/N��}bt��#8���k��T&����9�Y�!H�oц�=bX&�$HpWV�Ur��Q���wN��J���$��
T(�����WG�0ܫ�L�8�ҁ��1N�5P�}�Z�p1)��cd�Y�pb%�����}�qF&>���00�!���ûf^
���}-�y�f��'!4#_s�,wmCG�t��%��?܄��h�K�42:)��A�d��� j�"�|"��s�j" ?��BXY�u�~��L�I�����)z4.�H�j��U���Cc=�}���F�(�G��rb1-�d�02Ì�j��L������T��� 3�RTJc�ͥI��X�F� 5ꯐ#7�dĒ� o�>��b��]G ���'��_$���tt˶���Y��|�ZmlAX�r��R��X�ح#�L���ħ#s�FJ�Xf|��?��V�p�'Ի��P�	��l�o/[��v��c���::0�Zԭ6��m(��I4��<L.���`�'�{��^O�.`E܅�긍R>''� -�b-&��aE;g]!=Q��3Ï2�U�a��Pu�������8�\�-��X�/o�O�4�Wv%!JPj!�L'�.C�PF�w���>�B�t���P5[��(��v�j�0;Tt�˝U�X�"s�<��*��v����iU�@�q-Lz{�b=MI=�����n����sd Z݅����.B��C�0	T^������&��M�X������)���`���[�ݏ�2s�5+����P�~|1F��N\��GTI<����~}���/��V� �0�_���:?�����S����4�ԁ��rzH�3g��f(�rt*E�E�4����Q���ʽ��iů� ��mp�(|�Ѽz��(����c���,�h�U6�)�TM�	;���V�t�2��0=�14hH�f!پ"�Ф����"F��>U��K�1�D%���/���oIQ��ylx�(�oϠf�)j�q��a�Հ=�.���dg���ð$��X͝�&b':�$����7J��{D��A~L�n���U��8��J�����Sg�ݭ�j�F�mA��1[/���O���y�!❡���I��UrMS��g����~��0y�2�>�CI��7�������E����sf�A�0{��W�l���d�&<�]����/�vC��DUCFX�N�N
B�7��Y��pth$�ݧ����Z����]������l�@�hj#0�qY��M��>޼��]P�m.���Ǳ��\j���{����O�"��.�>KC˰��9P���A���b�2�f>�wy�5ս�0�}v�v�j��3�2��d#�<j�b�P��"���-T��n#S�Eh�[��֋���К�;g��&߭�w�k�������3��i,�Iw��3����K|��E�
�{���P�,�v��tV�Q�q|��ĺ1�Z�@E���+�`��hDƓ�r}� M�i?#8�N�,.�6��W8s�M
��t��K��\��j2�cV��6z��n��R����|W�/ߣ� #�f^���=3j�l�� t�`Jz�st+6�7�1~G��帹.~��*�t���u�mz�b�� >���Y-}�������"UY������}�����,��U���I㊬�ޟ�����t����d�Kyr�}��T`y�����<�Z"�ጁ&H�o��q$\��o�vX�[�ڵ�ӶS�6����\mq�,�%���rQU̮��1�j 2���P1�$�8()���>]���xg�gg�D�]|������@"E{�B��cB74�����Q���.�l�k�3���ka� �0Ĳ��#���6�?����	�+V`���5U#��O��<b&"�AR�7�׶;�0Z�O@�͊�o5�Fg��>N�&R��YA��|���2�/�v���2���n�4��~����@�ي]^���a:`���u��`_p������+�� ���NV�,[��H���Y���Zs;0�A�t��)���CX�VƃA�}]��e=���1��.pz�&GSH����D6�3i �A��Ϸ��:%�r�d`�+���$����N�Cf����o܄a�<�K�d��J���#ک�^�'��@ⱄԮɲ���D�C;A�bs��y�3����ƒ���<�g�e�&R�3��=��җ	�'�ѝXQ���?Ӻ��3,���������ꢇV5���v��[��y�q��=|p�U1m��BHj������ j[��
�%�0U��ר=Q�tT�X�<m�$��rU���0�M� �D��.�6P}�ˊ�IKK�C��a\&�cwf��V�M���l:�'��(5��	���>�|��Y��P��7��	,� ��5a�<	��jӾ������!_h`<}ef�����S�_f���"�����ػ.�����Z��#��Pz*�����b��j9�0꽐������w�5���h޲x%$ț.���
f�,]Ǵ\�����Xv���#�'4��Pݑork�-l��i��>����׉�#�TbF�6Հ�5v�J6@��G���Ex޺�f�j�O4��d���)�D����F������[�����k'������<���v�j�ZsN+��aܩoi��3..���"�B^&��u��'�-[��!�#* ]��S��pbӉ�m�����'5��	�I����·V-S5SV��.IhѾA]t���a��.��w����]-�g�WZ,%�~�®.*�M�kN�e�B�c�Ф�HI=]�f��f�Hݬ��wɘ\�?�׭����������C)ՑX��*��#�������4,�/���%�I�hF8]KB�"2M����Ҕ��O=,93���l�5����kRֻq�cBYtw��8�"A:� װP�A��vn�#&��4�����l4=��N�9�d-S�f0m8|ۄ��.=Y��)+v��9���sS�q����R[��9��^�*W�L
���Ѥ��5��%�DK�Qj<�~�~�9�zD�E���1�L�ԲWm�gs�T���9/�M<���M�f��5�<�7$�T�v�\�W��F}�$�����QM����C4!�%�����o��~���0-�8�&�t�m�:��~�_i�[�+�x�-ԅA�� %�+|�8���9M{���4��Vǈ@�|e���Y���W��|y�;<�@M������ZV�����l7R�P��g<��\w0 `j8�X��D�ؕ/H�O�M�����:��f�[+u� �i͊l ��Q,�G&%k��;������W6c*�I1r���WK�_�9�z�i>�Q�[���o�/{�҄���!�B�r�֍4�����"����	�=E ų��S�H��JwC��������K4�9�e����f��C����Q�x��ҌH��<�v�ӒuB�: �uc\�s��:�u�'��Q��AFU%���Z���1�;�so��HYs���M�-/
��l�8�g�1˶����}A��	�P��֋\P���<�4:��'	�z�Op�L�p����@�B�ts N_q�
�a�/cW%c��XI/0��K"F��t���i��rjd��"�;��p�Zn-1��*E�b:���.��9��b�=���Һ���9��g`˗���s,��o��u
=5ǿ�~R]��WRw���E�RE_/��\\T��@B�b/�ʅ�R�zD��j��6V�L��%-`�	����!�X�B-Z�T~f�ݵ�r���A�a��������Pd�6����y�l0��$БFhL���Sl��H�;מ+�[$֞b�iJ4�I{�#�3!B�(��2�k�j�_.�#���Ü��j s�*~��>�qHSe|,32��Z����u��)C{�޳�(�v҆��N���ifc�7����h2rm�Z́�!�X�w~>U�������|��/W�,v3d2j�+�E54o״�����í���`s�b6�'�n{�3!Z+MY�M4�e�����i�#��״��b~t6H�f~�K�$�9�n��������0������ƾQ�o|M���&yڛ~�qP��yzP�k1���b�B2E�1�j���Ia�@���;_���&^q#��J����H˘���A��T1P`���_������k����\2
�V<y|aK�&Q8m��V����c8�\�f��"��!�Mt�(3��`��]�0���bG9;���o�Ť|���5�o�kZ=�� L'��rjD��-�Е{['zfS�#����;��E��#��X�_��#��_�fý�����W�?A�b��̇k�ײ*�����5F���99,ll�U('��<K� �.�M��x���L�黈�b/g�Q����$e���J�@��H��][u��̯�U͋��	A:���#Ȓf�K얢ՙ�����ͮ��Y�^���������H�6��J-%�����8����؊�����-_�ȟ3�Ϻ(��ޭ)��Qᑴ�T�g�cN���AsS��گ~� ~.ˎ��3����]�8�&l�q+^�Ju$��\'��E�V���%j���J����=��I��DDh��>��"�Z?Ї�<��*E�5��Twck�����~~.���NP���� �'s�� �X4l�؆cex�Ҕ��� j8&�l}ʲ���K��Xl�|��.@���,�BQ��t�:'ن��՚�4Lu����Q�n�>��x���Kȼi�记,���ɫ<7�*�yU���V������4g.�՞��J	�8H����^�X���Ћ�Y��h�y��_I ض������{�Lq�.M��H/�~��4v�+�t�4lhi8���Բ�ZV��(h=���p�G� 3Q^�6�Gu�ъ}���dE���㳷�tx�ϥ:&q}�4����:�j����(B�ѲUF�j�3STc.�0��k������c���~�(���:����YI[�++=f�D����^�v�+')�\�+��W���>��VEXI���'Cy�����[��	d�cM^���g�q֕�Q��>̀���w@�z_Sk�ΟԐV(�u����=�tT���6 �A�1�Q�L�8
U���� �߄b���p��l�������
(=�~|��N�)��s�ٿf��5��x�cu�/Œ���tܸ��Fӫ;���2�C�=�����v���}�wU�!;i��U}�۾R�ent�W���H���A�"��� k��lfF..[p��@ˡ's�0۩l�� ���֛5�g �do�V��|Gj�$C�l�K]���	.C����F?��h{�r?F�&ʖ	v�aqK�uB������6��15Ռ",�ң�Q �W��[�y 'A���&���O�p ���o�O��ڱ�s�?pv;�0��=�M�R'�"�j(Ov}[�r����]Z�賗|Y�"�d.�k�b��G��a�:oL��~�4��b"����|�S�KSwPǕ�P��z^p@���Zm�tz�)�w�(�����4q��'�`��GF�|��5c�!(
<;b��lP΂Tq��^���x�x�j(D�.s�6ngŝԝ.e��t}ݼ�9'!��I�U!�T��xn�<�jn#�~x��$�	+|�P�	dh�B�}�~7������9ڛ[����~^�	!�;���Ü�_�\_oc�Q��.���N�`]�@���#�Ԫڭ���4��0 3��K�_�E⮞�(:��F�q3LZ(����R�L�%�f	�K��xމ��:}��Oy����S�D�3?1+��������1�{��[b���_�|kU����39�Wl��)����ԁ.Z&�Z<�c18;�j[g�@z���X���5J�-�[��P}4G��
�u�÷rt��`�y@�#����9G2ǢZˣ�S��꼆V���.W������`W�s�0�+0���e0ڇ@b��#�-G���P��n�PGX�u���@K�Ȝ�o-i�¾D(EM�1����?ǐ��O��2[`
�Й+@����{Y	�kZ+��<#j�lï�q��T
h���茓|�I@�B��g1%��A�d��N��Mx,����,�7������Έ �*�����V��$Ǹ7o�����K���@d��O1nR���K|o���/�xc�B�4ntЩ�31��S��i#G��#�h$I�{��
ǃ�n���d�-��V�h٧q����/>�h8��,gĜ��o�GV� �7~�1��C��0��:����W�usʟ�����Q�J���`X.^�ᣕ튫�+#�E����?�TÚ�V����x�[^��\ێ�"��f=ID��:� �|�����D�fi�N7��x��#�8���(%��V��J����7e��ԺZ���nE�\���賵��2�������Uq�	wK:��DҚ�kD/l�c�p	�B*L��C7�K|��c~��W�:����>�HQN�{�ݴ�Xq"�!�X;��<�]hJcC�ͳtH������˝gf��CH����9&zxc�il�_O8Ɲ�#Bm�6���O����1�]9(���l�ώ'12�@P|����ڥ#��>��	�Qi�2�,�`g+�D�"���i<ö	�f�<3i�����a��S�b֦NC���a3�+S<X�EQ�|��R.j:��9D�H��H�DS�x6�(�WR,{p`����ľ%d[�<��������Ң�=�v�ZS"�?5�����IK� +�L�\�GY�T.S��P�I.���vd�I}!���O͂%�28c"�JAe���*����:!!��h�֒㒗5%x���j�VEe選Y����]�D��A^�Hs��.��E�*�T���Mq?a����gb�%�DD���߰�Jn�M5��y���{Z�[Q���S�n*g��]
;�lxV����m#\� }>�hj��34g2�5���kZ�(�@X1�|���u�LB��vO�ͳ���� �g1n��R�*����7o:��m��Gs�rĎ}�[?�{��ʛIò)qe��Т%�0�@,�6�A>_�i䵯���ʱ�����!M|������}����r���8P��/��|�s�Uq9�JQ>��L-Ҿ>�P}du/\��~�g�n���X,�kl2C����Γ�t�����'���� f�M%2[�%��j/2�0�o���)f�W!vi�b��� ���	jQ�^R8h��h򉴧���S*���u$��,������'x�� �� ���hK����y.��m%��n�����/j3���n�]E&Ն�ׁ�KN��W��МIq��Fν�*�9J(��}�����kkT��L���Σ �òw�a���iǥfN��]���<�c���5�?��y�V�8(���.*>I�Yj�r8�ڳoֵxwג%e;-p�l&X������Mz�؁Xf����2���J��<�ϦR�mG���[G1�s��$��m��~�g	��(ȘJ	��)7���}~m:������ݷ鱍���������S��օ����n�y�P��%|�_����+�9O�k�Y#_n˸�mM�Fm���J��;��)X��J�v�e�&�S�ąخ��puܦ�^�%�N�Z��R�n'�c�T'��
�����F����M�����X�W�L�"/[jBT�MU[�0q�`��@#Bʲ�ۨƴ3�\�9��Δ�
�2n���<d
����PT%gp�j<M"��_m�s�sz8)0D��
�R�%I~'��H_�[_�u���A,�#3�įJ��x�<�������A?��B}��Nyܕz��9��2@3�%3ʌ�C31�� ��Wf)�v8See���:�Mp�!N^F���w��;�����+�!f��`B�3���h>��N����@Zm&�ܨ��t}%�R��i)6÷x=��Ԝ5/�z�*�A�����~�C+8ļ.{����"�W��#M��2p�bAӲ�!Xz�ր�\*�1�/t"����A��惦)/] ~v"O]��2zH�3�*:�zw���7Ba�B[9�Y��Pj��֐p�����Cnٞ��զ.j��:n���
�2sS��cs
�:�`K���V�e�;��,�/�>�_�����ӣ��|
��{�B�G��7�5��uoݮO����ҴhqT0;Q�-%��!�שׂ�t�λ�%t���Ҹ-)�'�`l�GW�w���I�+t�1�+7���Nu=1!:Y`�p�l��f@�ZUy�nC�k�b�oPO�`7���x�D�}扻]l{���sՇ�7ò��\�E�Z���xW������;<o��S��R���Y�ޔh����s� �k����V�ڞ�z��'T�+�]ί�XE��HR�|PpU�r� =����o0k����ׁ̍����c�`)n�<ڴ��ģx�j���<�X���L����yY��Tǆ�3�{"ba����"���^��v;1�i�
/K�'��D?����0�\�,�4�fk4�qH���aJ&�������>/l�xk�1�|<tEA�����iQ������� ��`��eSyO(���	��LO��C
4�uDȲ��U���ĕT/��)�/A6=�v�ڻ��:8���;���a�� �Ǜ�o��Ef�����j�V��c�O���d� �q]p��p��DOTtǓ�ʞ,��CkU��Nd���� ���CXnY
.����/�����\�D���~�J^�f]����D#����/�(#1m|X�u�x�a���k���	T�m��B�SP�T}hjc�C{!�9Y��P8�"^�N�p-XMϴ����9��&��B̷���0a���U�h��.�� =)�YA�HXW)� H9(�m�a�qE��4Ok�rz5�r|=?����r����ԭ�p�ٶ�i�EbW3���l�ˇ�]a� V�M�lU�����@����.=�y�-�K��V=Iy�����C)[�߰Fpc;�+�k�����ż�:Π��>��������u�RX��S�Tv���(�^�O^�������	鲚������L�D����ɴ�X�!R��X<Ա��چ�ͪ ����zc�C]�W'���f�bn�O��/�^.P�{�!]�<�i�(��x@��w G�����[�b�M���� bD?��Yz��%�F?���hn��g̓�ӱ]N�uR�H�SRYqJ�K=�>���7�0��������=l�bD�C)X�o��� �H��V����t���3��;��j^�BC���g>��~�fm��i/�����Bk�7�p7C�����:`�_�ɗ�Kѓ�;0��П��2[�x8��D��0uo�iMs?Kw���%�4w�Ѩv7i��X���f�g�S�Vԗ�S��gE�f���i�W3A�@�p�}[<�5Ӟ�#�F���.�A'§�ye�EP����~*��$�8b3�07��a�A.*���-��Z�'�X�:e�r�!�		�;r�P]bX��'��P�R�5D=vX�vx2�_�*�ѷ�G⿇��
:/Э��^�*D�vU�0��d�+�I�	uZ�m�C�eT�r �jDN����à�i��_�[="�:��7��K$�E��(��a�Z�&�������K�3<+����k{����`�{2nkfKE-h�5�]��;��u���ԕd�gń+T�">H�@��\��A����x������2�Af5���T���5���vl�����ޟ)��Z��M�w�-M����}�ں����1� F���̥�.w���.�5�(�G�����t��e����mA��QOHu@�������bpX��Jگڪr�:]� �/,v'�Ӊp�.w*ͼRyC�]E�5��L"n�n�
#�ť��W�(��w��n'�����M7�(��p�}e8q�ڼ�{�L���)^�ľ�Ȼ!&�*��q�9�5��,� Oh�r����undky���F=�˽�+Q+�(vVx�9�>~�ZVG�x[�Y��͂`A��w�|�L;~A-¶��Aw�s)�?b��A}.�n9B��v�n�wxXE@ l	u2n�U�<��lh��7i��O�%hy���\tӻR��ʧ��T�n'�uQN
P~-��oT�+]���j�B�����tt�Qy��S`��e�L��$$�w�����k8��߂�K�V�z���wӍ��m�]��7��+=��s(�lR5��0�?u[��E�q%c��Z)C���/�m���(�{} ��%�9��@�^���%�}x�
F*��6ߐJ�i���R��!���Ò1b�D���ˎiy�6h$5M�z>�����ڜ�!��������/QD��q��� ��D9W�
��$�﷗��1ϯ]�Κh�r���d���|��9ڋ�t5�t�F/��X��02%�W?&�q��t��i-�ڽ�%�2�K*-ɹ��eW�v 3IQuu:��qʤ����n�L6r�z�J=#[�r�nїF�3�5�(?lgH�t����.��>� 8⃼�}$�iv���E������^�7�S�����@�Γ�l��ڡ�?(�OP2�t+w�aQ�ή���zS�#�Y>���U���i����5���3+�}MGB����X��s��-K�S�\����I�97�|e��ӞS%^q��lp����]#`�I������O��E�<�ء? �'�d����CO�c�=��win��X��~\�ٟt�\�)9�c��Z,���0xo	��Wޭ��;�p=X�M�訮�V���g��縃rⶢ�
���z���RWTdH䡣�IK�q�H�-�E,�J�vg��I�0�����:����08S��RB��ʅ���e�X~x���q »3���q`�y;�Ko�w���v�����6M}�HU�Ά����O�g�=m)��֮Y��+��t����i�禍Ԡ�E!u��2�������/|"Z���A��I����7�C�b�j蠋f���B�7ۙ*y����J���M
�f&�|�ۃ�>�O����		�#�`օ�xr�:`7lx���'nR�H1�)���A�]�ԾB�����R��֛9B{�Ь>�>�Q*�v5�O5�!o���� ���t������'���Ss����R,s�	�|������1]�?G��{�>��k�����Ęk������J�$����T�_~^�{�
�$�{W�d_ɿ�3:ED,	)�R�;*�ǯ��g����P!t�4!��g'�!�F���Reh���3�S�P��lO݃ ���#SD��g�&���B�������4�[�4_�WM�2x~˵c*��:?r񲹴w������ pP��DyT��pb��e4]%_+sCc�y.��3J�w�i+�}P���5�k�~�"��WIy�ֲx	3�ɂ��;��hR���x�:c��Q]\�� ���OV�3;��g[�3�����Ճ�����9�ڒ�k?��Yg��v�����c4_�ג������C5�7����ށ�?���s���%$�t�F_X�}A]�g.aD&Sm�.��,�'�FU�M�q�UwIК�G� 4�sf��\��+e���
��5���t���Q0��Se4�7����?@U�4���5nh����Ig�Ġ��ك⏄"�~t9AM���b$�ػ����:jfk�s'�;�A��*�cRw�j��L��a4^��h�I�Q��[�8*�;���UA�Z��)�ힿC���MͿ��"��@���p{X@uO��=��)���*߉���]����2<� �E�H�q�cN� ���w?#B��J�j�t��v�L�*�B��y�j)�f"(�\߯Wm[>�k�f�x*�4�6��4�16DB��NS��h�&���[������c���c��i���:ڡ��}���`gۙfQ��L�gW����5�tx�[Qvu{�$���{��:���H���t"�I��V��Nd����H�k$m+~�/�aM�;Kd�ǪXb���
���z���E�4/�&L��d����v�_y���O}����/���([w#]ŕ�����������a�O�� ���8�'��phO�rJꮭs�ď���r��ݪX�7�3#?3i�;t">�M�m��e��6�gk�vK���&��,2��83Ŗ)7���8̴�����O�2Lɤ�'(;U��)0�T��f �T˦�P:A<d��O��}N�`~"0ש����{TR����|��oBx5�J��ʋ����/ڬ�	�i%��P��֨L[�r�B� ��龬&��p�L���_.P��͎���Y$xK������^�nv�B��S@-:A��V�XXph��/��f_5�V��6:�e
]�n�+U��K_W_x䵖�R���ڜ��e4n�%�Ѓqw��R�ˆ
�"M�xZ�jX�L��<'�3��EBW�N�n��?��*:ZM���u5wNc�R$_�MG1즈�����:n.��xl_pB�����g�|O��p�?����l:�1����KI��˫��5o�̘G������^ۋJ��Qg�6�������}�E�h'�b�	3y�����G�t�j�xd�E���g@�Ӱ��ب�mϺ�m|L3������֫|s���~����ᆥ�bꚱ���8-j�Sz Yɍ���U�ç��jV�B�ńu&u���]F?�E_>Z�I� 
�]J��DzȾ3+�lbW�}�>�]{�j�on2ͭ�!M����s�tL����#���N�����5��p؝�bnp�{!6�-˄k;��W�A	��7(�*����mj9 �yp���a<Z������'�o��܋�v�Ɏ<J��(��w��Q�?�����R^1���7���}�Pc�>�}�\��㗁h0\<���~݄�ѻ�X\(��uh�s6���?�{����ʳ�F$�i'��D6h1s���,�=@��gΞA�K�e�1��A�� !&^˜M���	L'�Agj�~c�LjQM���_8��Ld��[���(��m�D�t
�/�B�{�(�^�b��
��伂˭f�U΢o���Q���y�^��i��u'Y��V��;�zzu����YPF	>��{���NC�"�i���@� �W�@H��Gv��E��
(��R: �)nR4���'�2�8}���fJg�̐����R�]�{��'��o���ڪ�˓���Ң�l���?H���i*��t��-j��W�I���Z��|ܗ���|��g��ƯDe��Tz�}��n����<�D������z@Nȅc�&-��^�D_�8�p����}��'`n�!�)[C��Zsϒ���i5��Y'� {>�Q'{��vN�+���A��&��2�n h�7�q�%S�mFq���m0��T�!���N佔�#"Z6h�l�\��VԞ������������r�O$~�`���"�k���p�4��)�>�_)`�s24 ���d������kc���c2�,9�9��ʽ&�mu��پF��*m��B�)Y��q��Έ�B��G+~/���Oe�,�R � ʀ]�(`�W���#p��L*�Vk�mH�|z�i�oH&C�L�I�1��O�e�{D���c�݁����.��'<��3A�a���`G������ʥK�MK�:E�9�|�~��L��Q�4�!(�W��=�ʂ~s�N�0i�c7>\آ���������e��[M�]+��-�Y�5�؛���h1G�o��Wd�i'��?�\ �ST�A�@���^�}��V�c��Y����!.5�TQŏ����a�%Ɣ���A�ƽ�p"<1Îզ��(�0Eek�7!\�W�od�Y�S9�˓ۗ�ǀX_	���Ɂ~fB4�
�&��<ˍ����7@���ߚ>o/>�M���]Rr��+�H��F\!#-��O�j�b��H��B�_Ɠs��z�ѥ�?�ZG<�NZ��qMY�����$3�7U�'ns5��@��cFy_�[Z�L��f�,a��X�٧K�bZ� �(>�Im��?��V��bh)PP =_�-��:��y�B�]�j��B��)$^�Į�k���\a����k(��l~���"�_���^�Π��3Z$�5�r�e��Z�q?�����?0Վ8��^��Gv� ;$���ɪSǛt��R�X#��PR/�K�+�6�	��!�I����FTǿY/��Tc��;=d�f=��B�;�ܴ���(?�Z1��I���R��տ�����s���p���5�\&�RA�:B�ݪ�LL7���|�<�є&�����܁޻"P��e8��`������G�����G�x?; �f�̝$�Q&Le�䨻6�����Q��as{�-���.�ٙ
gfN=9? S&q*��ŉui=V�*�28hd �ZÐUpu������I	;9+�sBXuQ�A=�Ç�j�(�.������JD.4�k�'V���>�X�CL�K��چ1A�̆7��G�a�q�I�����Zf��i�>,E�����	���C�5�B�E��۱);Q)1吼Q0�6`��\v5����L�E|�]�z���Q���M&���d���
��L/����Q=������9��v��,GFM��Q��_�|!�����UB2J�t멷���Ds���HU}�?��1�	{KUYR�!���z����"�<�� �Y��&逜*��� �Y@��
GZ��ZS�Gx<v:�+��7� �N�R�=��CB	�����.v!L]��t����Q��(JΒ��ɖP�S�|H��}�D�ҒX&��[��u�×�j��S�z��q����g
���v�F��F���� W�@BV>LP��M�k�7�O������s�c%��PB�����ŽA�v�����p<�w��Y�v��\��X��ez��K�� ��07>�s�/4uB�vל4�X'�p�GA0*��'�����p{��$뉤x|_��Τ�ۡ��~�xY�����h k��k2W��V��Mް��JH��Y����YL�H�i~C:�4Q�� 5ݫ�|��otگ"�WF0��wi���:�I�Ԃ�N�v��W�7(����x�b?�d\�#�q��4��gh$�4Bbg�OB���M>�|C�V,�`Ulx�'�Ň�'f��)��#��.�D��c�E*l��~��g\E?���dM���ve��x6H��j�[������"����m�$�]͠���6�׉��lV8aƔr�7I��F��{�.�+�� �z�A.�Y���g�sG�%��WӪ�4�l\�s��Q��
�
�
�Â�kN�Z��0�IB!�a��Sy*�ʠ*D�N�-5W>T9|���dl&Չ�f�\in7i��A�G�OZ?��GOۭ#G��C	��Viq_�J�������r��+H4����k���xᗍ]bDP���rj�^��o�/΅�C���� y�-R�Ċl-�~oL������npe��_�'��@�ʝ!�C��sj�����˾TL�ʅ��P_�%}>�ѵ&�- 	��	Q.*��D@
������+EjRV��)L�-����T�NU��ma�,���-ӹ�+`[#��-�O[�����8�-x,>��l'l��W4�7GQN�8��w�\�- ��2#r�U���~������T��ǍI��_~)sq *jl) ��nR�^���턫�_�'��dC��~���>�^6���}O�������
�fs��Yx�J�Ԟa����t4XY�+]MԦ\��c_��y��f];���g��Uv�K��~C6�)�9���6>s"�����U���HA)���=o��Np�)ɀ�~f�5w�B|��H���n��F�j�����.O'� 7���yPgV��w%Y�%�S&�@R!�Ch6���/x��-�`�ئpR3]^�(5s �׋/�w�%D�������-�-PY��1f�UCy}�7�[CL�Hs8��[=�mY�	��NwD����>/�45�;`�n;$fm�����c�d�Q�uL��ʴ��Sl���B9�EK���l�����b�6ˠ$u�
c����-f��mi�l�a��Z���q�ke�ȫ`h��(/������ڼu�҄����ؘ-SQm�!�+=)ܓ�t�'R�%�i�@��k\�A@]��^�J�Wl�s�h���M/��-���I���"��#�à |��=z�^sz�}H�1z=HX8��t��6��6��Xzne�+�Z�\.+� �Yb��N'�SB����Z+E��#؛��m\��A���OO� ok}�{N{h/���"Zp��_�L>��T��ް�\���� ��#%zB���F˒`��p��͈�|�/W���#�n�xs�S�c�G̥��þJt4��_W�ti�q���s��/��K���}�躸T{�5� ��x�S��)cR�A]�t���)Z�n훼:;\��:��h��?���u�g���s�[!mm�����I�߼�M�205�cp˅������'�fiҤ�z�ЗyzD"b�|.�񌧴O��w�$�0��ލ?��@0�֨�A�B�+��?{|��W�XOYC"t�~�[��Iq0&�
�=���e���%��=�<��[M�]����F8�vJ��EPw�(��x(S�	��&:�a�sm�O3�}��_}6�@qI�3�xd��l�i���O�y��6>�:���( h��|ρ�����r�R�'o��^3v�SDq�E���$$�MI�Ԩ�[胒֪� �/��ˇ�I���AKK��9ש��ɍ(��;D���*8�ƎOFr;S�O�8�5��}s�XhC�ݑ��e�x���yj�o��=Ŀ����.�A�˥Mw������\6���(X��������
�Z�@d��y��3`n-��ܡ������8�oҗ�zY.���%�{���+�wIr�9yȑ�O����*菞���s��Z�=4�tH�0 g��h�c0�[���j�4�pOn�y Gb�;�G��NP�ݴ?ƒ`�V�;M�aP$|r����x�!�{Tdn���|.�����ڀK��5G�F4��> bsL����v����UHl�� �0
�l���d�/��6���Y�$،��Q/�q�4�q����.7�P)ٺ���o�
3c��-���83܄*O�"r8{v-j"��zp��/O�Y�7˖T���f��zw���/b97���������Ww�������u�c�����B%o@k�xtǡ���` ���ml+��R���_����VY�}-���X��R��ޖpOU��ǹ�g���e����2|��Cb_�g{՗������t8���SXd�h0I��#P	LN38�yu5��ɖ�`<A�}��c��zq%�MkN����c2��r%_�����<d5�@¾9Bl`���$�' �_�^|ƀ�y�4=�;�.�	̀i���d�9�#sG�|��  �9�Hg�>N��#F-�8�9�����ų̀"XJK�mbU9��`��V3	DY���p7AM��?3(lyn̫��6c�M	��t�kбqoIrx�|��D���W�H�����1����/�t�i�/�%��#��(}�o|��?���w�^�rK�UF�f�n�~ )GHM*i�$ab���p�^�ϧ'�β���DVq���ra,������̶CQZ4ΥV]^!���ի��<o#ttt3����Fp���3� � ӷ���+�(�مŝm�!+�$^솒�pE���0�J�Tn��!���[����;�	N*Lm�d�>�w���%Z\o��<��r��<c�p�H����˵z�_	�S�Yݘ�m톜�X�N�l�<�ޠ̴z���y(�V�١����_+���!�B�M�P�\[����px=�e䶊�� �jk��T�V(�w�%��~��Tu����?ۍ�߮:c?�f�v�@�]�$��\cYj��yt��;��w�!*�j�V:>>� ��*t0N���̨?4���S�Hʵ��: z��!�^85@\'���
{z�ѹTM��E���$��9k��}k��;���SS�z㌦$�1���4�Ьh���� E�Pu���RX�<7��#������'���z�}���"�B ^ؓ�Ϯ���Q7��˹�3��.}#�I���j�j�Z�9Y9��%Z�����]�\�,�caCg��oF�|�B(ӒZ��=�����)=�,$�]C�iR$�z�5��\#/��ĕ�ni�����@(y3���w��� Y}��/��ޥ��ٻ�?�Zd
��6�G.��I傕���ᛢ����G��17T%��\^:��u���i�f@m�~?�����`��Wh7 �aa���a�U4;�\ 1�&1fjNu_�R���b
�̢�Do)��Y�a�K�d��'�YQɬ������o���J����[�1ł��3K�ԋ� ��<آ�vwq�o�U�j'eJM��EJ{3'��üڑe��yta��m�w�J ��7�$�r?���hOLvX�������}2{dz���a��<*TrH=�Wŗ��6D�'j#����:�  Qr���Ֆ�)���|��Qˠ��JO�F,<`IH����N�����gK|��UNYn8�M*�_Jv��O��j�f�������^
�Q��X�����9��}�����y0�DO���º�+>����I?M%�Q����{�E�˹-�a�l��.�xa�Ӂ�
{+���\s�E	���8�{�����?:
,���%<VR_Mw�O|ԅ���&��2.P��2��O�����x�+@e��J�ʚ0S+���ŢX@J/���h�����3�NP<f��d�����Ֆ����eL޽�H�RO��*���c��Mt�Z�Yc�XW��2ށ����)Ds������GP�����{g��Q���!���#j3H b1����'���L�����TOՓ�?�C-�fZQ6��֤��/[��}n-���\U�&a߻�f&�^��.uĽ��MI�)�,�.�k�Q-{��t�c?�� �^�^BG3��O�T��C�,�K��_�Qn�,���wЀ �����vܛU�q*ޙt�����`�K��)s.g��D�-s2-�Fi�Fp�d-�x�p)�����jQĜ��StNǄv���D�)Gk�lI��$&q忋��p*�IX9�w7Z�4���l��&���-�� �b���'B��)V6�ag��u]��g��Ꞻ>Df:��f�c����by�E�{YH�qs:ͱ�`v�fi����b13Hz'����`��p~�j4S�j���G��2��s�2�]	=k+�Y�qX���{����F��<��#W��:��6���O�cw� ă?��D��*)�"�t+�xl����oc���)(U'D`.v�m�>QZ�{h��"���9{���� ��h�Z����s*6�}6�����&���9�
�0�"dlB����6�$r���T-�(c �V��-�(�	#{�Bҍ�=�"�������~v#�����})79
�<OX�c��"J��N}-���(t.֑��gڊ.T`�>��>�]ah��MK��uD���.N@/�a{�9Z	��U�۲��m̈5�ū��ĝ��	�"yM�I���FF��6�EX�1L�Y�ɭ7G�����^�d+�E$���/'F���L؃��G͋�m#��b��|.�Q�'�M��t�q����D<���
sN[���Q;�d˨�d�]e���[��1��|{�Gъj���`Od.�vas0Q�n>�c�	EO���'}�pg#�.�v��F3Ҝ�����J��i�?ni�<˛�d��i����SH ��K����x#i�p������5�[wQŇ#2��h/^JS�|���otk�z�}���L�$��]���eRG�U�E��}��5ʴ�¾X�j0��)l�����3ڹ��Þ�����z��'0/��J̮dU���-]#��nl$ak�D�lx�|e��;��ԙZE��/o�{Dc�z�a�^�1��K�Wթ;�>Cp�T���lQV�R��S��?2LAn�{�r��vD)~��*!�p���>x}L|��}7���2PɆ�ՊX�,�e{�.��ϻ��Ǐєhh��%e���4ྙ)��]fA�Z���'6�����זi�EH�*X�x���r�Y��s�I�Y�!P�z�=�q��o+s�:�=ৱ�2L�w�A��8fk�oU�91%�uo�X�}[��MZ��� ��i��Y��X׵}D�����r��$`�6�?�hGNʇ���L9��|�lV��pJ$��e��NL��^���m	�ӗ�z4�t��֠�f���3�H�+��;���9�72x[�G�e��G��H��{���\�Z�*�`����2D��	w����$l�et�AB���H��鸭�ϯK���h�����RZm|����UL�j ����v��60�H��a�'.��m��`�% ǮI��ƽ��(g�+'���u� xۭ��U8�--��k��7Z��4��6�%���t�$�c_޺!���Ѓ`H����d�Ƌ��Ӊb�f+/#_C�f�\.�ak_eiP.ma�|�m|?�� ����0*��W�z,�׺��5�H([E�|��d��,��`��d+En��kBT�+G�D��Z�� �*�LJD#S�1�(�6:���\okz`�:�2KS�K7��L#ψ�2�x�/�a�5��n�X�<�?����|@s���Y�Yzl܂�(�b�G?��e��u�*A���,tp>L�ӎ���q�I�43��q
KN�
d&�8�ʋ�x_�	ol>1u�u@�3�]�*lQ��I��8�P7�]��6��hn��&�F�h^j���[ɹ�̦ʿ�Ö�8J�}��,�~��/������hG�}�T��7*��q�@E���J���濍sr��6�ç�mك|���)Y��N��9��b��QI��帄�6ȸ �(���jٞ�n�[�ơ����b��g��P�`b�C�t4��-(B���W4��A�\��#����,�]^aB�����5� <�;cy��&�3�a
2v+�T��F���Bk�x:i�9�4b�ƣ��K#�e��iH�)r��ũMh�qn����pE�:O.q�K�O�;�1����tzj!pp�(�ٺR��'��~V���i]a���*���9�����֚.��rkNbF�v�K��ȇ��uҝRqÞ�A�Ey�kn��
���>�h�h�"�Y���v��������@��㮦(���"�.+�s��AFmcj�J�/������F�|gP�`|��{R��ʑ�'�2�Hmn�{~;�U�}�b8�� ���O}[|2~e�.�|��zϤ0𤞡�A!e��ci�Ll����~@�r�Y�V�)��B�c[oˉ�O�O���3Xd�q�,��g�^
]�(��d�{�d�1���}�A�����3���z���E���X�"֭W;V��`�{�?,�b�(�:.����X~�9�u�D�'��\e���֔>E[3����N)Z��������9�ł�P�½R���;��vK��w�&9����^��j���J��3�ou�xj��q�A�ˇ�Հ�,��"(�/�������֡����jɧo�c0V��}�ޛ�g�<T�`�@�By1h���Z/�S��M�e�3w1�z�-ٿAy(vH�6I�z�y��©�Fگ��3��Ԛ�o���*W[C����fERO0���C�Bȵys;�0Ž��3�>]n�J�nðy��ǐ��6ȅ�|!�����$�su?��mOI�W-y��������El�\���C�М���Ю��Y�]�ȝ�rg�l�{G�!u�bÎw��I��	U.���L6�TfF,C[q�V�z^n`����S���إX�2�ZN�[A��̓�z(r�|�@����t��'�Oo������ң+�*�c��6����K�Kfw��>�1�7���@�>�Kʞy��ʧ0�/�<�Ք� �qc�t��I4̀��Rf1m�'��=tJ�顆�Ƌ�䆇�a�v7]��SE�]ql��6s�%�U�>�U�2P$����_�#�E��NĀ2W���u4��o��:se1��u2B�t=�AH�E\�|�����$���ϕ�j��i�]����c�++��l�ΰ�L�g�I���1o�<m�>�9c)��M�)s�辳�|;�͚�qH(e��)F�MFACP��ո�Z�}sE�� ��Q@>+T��'z.�q`�� �[^�;�B֯�%�a���!l6��o����>>���E���X�p�+�\���o���HXn
�����e@���K��B�����~y(�h|��4�,��D�3��w	�[F��F��� ��0��(	Z�<�>���g��Q���u���Y��qm�Ѳ�,r_%����o��l�Z29/�'�hi����aր)�z�bM4>��U��L/�$��BI'�=	��P����DlX���{[V���C�0��d^�Viu�#]ͳ�6��h���	>%�<�>�����RX؅���#���{��k$��_:� +��
�u��_�k��Rܿ|�ѩ&ћn:
]w�E�N�6��2�������o�[w���q��Jz�2����?z%B
��#���:B�s���$^c�j�}@��]�<���.���]���z�a�����^�(��Hz~�̦NDS�7�ېuX��
E�Aƕ�m�4�3ҝ4'�3����6�����:�����f-��Z��1�z
��8v���W.���H{G�%���/���검��ԇ�}��=��Ɔ�,�w��*�f���a��F;���!����#�%mr��x~���n4.��b�d#���8-V�f誎��Ƚ���]�ȓ\������:W>gY4}�E���n���C��#��[q��A���������3b�>k��)���D�X�'���:�r��C�\�,��=w70��1w��9�'�=�ɜ�A��$[^�ckL��Z:w���l�C�8+���ӷ���#��*^'��p�gS�Hڷ/e�k���T5eC⡽q(Z����V��n
GP�����Yv L��"d��t��n��lE�R��(���/�x$�Ѫ�e5�5{����*�Q:f�q=u4��2wQ��D�Q/�u���&k�?��:�3�K>Kc��-�W�g5���4�ыkȚ`��VN������&�������{�b��ΐ���?�7̛�ۉ`|��_sMN��,W 琏�y�5d(-�\l���;vQ?�䡽pGJ����0���y�t��:D��e��IO�+�E�4��]l�Q �J�N=>���>"U��Kl8���5����0X���GF��]�^��CN��&L�8L�W٢�?�z�H/����[&��AV��Hv�G�n�U4s=b�����`_^)9r�s��p��mE��$��Y�gmF/Ug�����O���܀E��_5@#�-��3z	�u5������LKc'�p
Syq5��9[���$���'{�\[��-���\��*�#�)� ks����G(��=Q�=2>�T$��^�̄l7ڛb7lg
��H�=�{а!�Tܽ���2�u���^%jΘ4���s�ߓ$]�,���b,D��]/A5������?�����G�a#�ZƷj�6������8�# À��%C�Q��rX������ϗ��j�=2�O%��#�� rDY;w�"u��#[�7�qvu�{��{���V��"� �Tl\6��m�qw1N�-�:�E�]��ls�Ǵ��u'&}P������z�R5-�&�]���Ns+,?&p>��/��������O/x��O'�|ZA���X��f��e�
�޲��
+mY�"�I�� oj��Ǳ�$i`�R�L5�;3�5�eJO����cL�V�- ��R��Q.b��� HU��
i��P���W��X#F��HN�SB�4
02��X��r�j3�'Õ�e��r��@�i̊�nm�UI�޴�g;2���׺�����<����6W���i�Vӛf���i���Ko�L��?q����EW�$}�A�z�W�J��%(�$��t�<�ɇ3s*��T/���
�>R�#^;J���fL.���Z�	�l܊�_i��=�E*Ք8r��#�?ˎ����?$�vi+�4�:�U���-��p��
C��v��˸�|�D$�����C9�q�� &c����41:��trO�n%�.9+�o|9�c�1��_6��UU|������xe����L]�c�m��e��d��M�.�!���S��Q�@� s�]:5�z�6�3
�� 'F�F\�m������E���}�r�f�a�� ~T�}̐�IV~�x�N'�� �{����c#-Ay G��rp�h���ԇ�I�{(�~����we�,�����S��sl4:�%�z�zV�)d�g�LaRdvK4��^S��k�	�ɇ������p�<�F/������'��ggH�,���*<�$)t$�u���R
�@���˥*�Mx�Ć�z̈́ӭS��g�A�_p|d����i+�T/����Q�B���f�U�0���s*���9=��/$`6��{t
$Y f�7�k�mT x$(a�
�T;�8aθ8��»�V�M8h���%.�5+?�r^������;���	
�%��.}���(gdys��3�n"h��ɟIB���ۦ�����|��d.�P_�:1A��L
Un��T\��)Ũec����&���)ޅ���B,b���� K��)�E��*����9d����2�~P�m��ې�/0���Z34�Q@�sh5�����w/��XO4���Ȭ�C���������u��̻d�����e��N�U�1j��)��a)��V
ӆ��L@�����)<~�J+���
���sʬ:�B-Si'����Y�ECoG��CӆMV��u��B(�LH�֫Z�d����z .���&�
�6l"�j�=�	d����f�o��kKl�n���%[I�&��e��Ku����YN���f2�}�6�p������Q�{����D�3a�؞��c�R/�ƞ�F��z6��c'�-e\R�h��ͱ���� �M���3����1��N���	_gO't�Y���>5�S�������L^3G��J�Q�m��X��&E�lG�
H�(H�YE�t�[.�P��� ���iՄ�
��gQ�/��1�y��ꏘ��<��nF��K%��>��������A�+�{,�Oʷ��7ڴ�0��3H^ʹi+�?)'�>�m�`���J�'n2�v��&�?��޻<.�3��~r���aRYB�#!�^.��(8	=ʰKJ��h�B��P>u<�P�� \�	c����ϭ 7 �u�yqJ��I��??C����`|lI^VֽE�����xR6�$=�a�ן��g8��]�-���Φ�t���nȯHU�zF�����L�i���j���rY�gN���^	��i�ҧ�B9�����e�l�0��
� %�J	�h	�)��><�j!;��T�g�h��°��.��*qp�Yp�|�3�2r�Y�={��G���B��˿E�!��9�B��R�۸��0��8D��v�@��e��s�	P���.~��O�@�k[��.��@\ ׵�.a��Cz>a`��5!�Oo�I�����w�WL����Z$1؂�p�I4}*3�(�/�dz"4�S����'�C4�&H��4�6��7d�Ӝ�G�j|���Al��@ E}AL��{Ӧ�s{#�[�����������kMڝERv��ׯY��R���Rns�� ��v�eE)_sĺI�A!�Z��1��5�
��%5Ę]kqNܟ:`��yL��3`��*�W�\��";��dI%9#��~��v��nt�v���{��܆�+7e�r���[q1JXW����h����%χ��3�A��С��EK�>��!7FӍd����m�a���
�"{۩�r;������iU.����u\ì���ڍ�tD �FN��ͽ�Z�.���"n�a�_��	�k!o/�7��{�� �O�꜉�}���ݑ�x{�F
�ZW8ly���E�aQ�����"A���|�����%O��1 &_E	��#�\	�o�+s<oxc�G���Z
�+ֿ�޵ڽj���v0|b?p�a��y��U�;m:�k�UE�ȸD��+��%�b�@R[8Eã�� Sz�{O�ϮHV�Y35 ܒ!��3�'}[�<IV�ЗWg#��������96bk41MQ���C���f%���l�B�g_�\������#H�D����$�3����)k"2:騸�7���'~�a<{���X&�׭���~��"�~=�OUR�vʹ�PZ?y9��;�[5톒%��h<%�*5�����J_A�Qz���}�����:�L���5���+>[&�� 屸�Vҋx�g�+����n�~���X���8P4H�b	8um�x_V�m���p�-���dq$��Rj�o���*,3LU�D�_�E?�XE ���"PGk1�����H�s�E$1$JL�g����`F��s�G�H�J�C&KK�� ��ģ�IЪY��l������p��Ʒ���yo䮆>��|� �-�w6�I�J���c$s�<g|6�D�O~1T3Zh2S���x Q0߫ڪ���h\G��h99��A�g��M���_e�6���EB�c����0@���n{8R_E�6p��A�g<�v��S���/���>�yٖ`54� 
��T
��������)�0S.�-*K��pSt�*�O��&H�9/h��k]Ӎ��ҁ���>���:F�!�+�����#�]�<����~r5B��2���/P�xhto���lj�P�4����I��<>�lǱ�p���k��z�O��J��,b�E�g�1�n��[)>3����+�dWf�����)��*ͭ~| M�(8�����_:Y!Jp�o���L],9D���1��\ɔ�j`v�QȤ�)p��� ���,eR�
[�V�<P��G�Vq��;]k�)̊짆~_%�rK�[ZY���(is36��7e�wy�g�"QbO"l�Ͷc�؟��ա^��s�w]���ӼN����j��ＧzP�����q��r(�t�.e�,B+$�aW������[΢��LR�4��$!K�Qo>�7�{�o�꟦跓?��u���÷M�o����_e�����$�k@��_����1�6����:S�|����Ϋ� ��vNk���o�eX��F��>��>Vy�|ЅOq-��$�����fk�诹����
9�ɟ	c�b>�յ�ʯQ�9{��.�LC�1�l�C�o�e��\���������8=`�n��l��77��3�U�R�A�s�Ӗ
�S��:��F�<�t��Yqx���S�Cr���&�HW{Κh�xn]ZV+iqNL6�`��uX���*�����l������Fqn<��?�!���1�q�}��s�ōv���?�5�qٜB���Z��o\�6^�(ǥ�f7��_*J�ԂU�r'��i.+\��׍ָ�W�zW�|c�&5o�j}�c2�Bdj��-�+Le��̒I���ب<0)��d?8��d�O�'ݽ�p�+4����85�p�t��CV�%W�ռ�˱��hTs�����
��̙w��{] 9�G7����zY�!�|ha<#�Tĩ�|��!��qU�[��ϙE��)��	����걨\�\);�b��adUWlYٱ��sQ��'�9e#���ߐ,Z�#�&�(��S�p���ox+��M����2���O�(��7/X~ �lDQ�j�)�.�ӫ/��46�%%E���>�x�H�Sy�.�m*/���Z�.'�{1�|*K&s���me���� ��g҄R�Bw�W�+c��t�z�Q;P�W�D��vV+�}�pb���rVʨv�>=��.�Q#5�g�������m$�2ޔ�+���a�����I�*���V���K7��6����p�� �?�M	�IdْQ�2)��T#Ep�\ھ?v��� dD�p1��y������$2wG ��V���	b�I�G5�)���;2�.�ߞ3C��G��Z�*|�ɑ�m~�ke�:��)�oЅ�J*:�k{6�!��	�d�Y��QvN�# ���=�O_�;,j��<�my��"�RIb���&�ڈ���*)�ϋ��$���9K�9�d�-jt�#	G>ϗ�AԤ�����]�ys�8�;7�9I�vw~�;Ǥ�l�D|,^M�(е�"ϳ�;Qv	�Ǐ^�ޛY"7��+�t|�3�V�^Q��;F1�#I:y ��lGR����j[6��=o�ż}
b%]o�a��Wf�C���E����-߱�� z�XN��#�����C�t��$ƻ2	"���)����Qte|v��~��GCf�^���u���-z�P$< &{���n+�C��aSi���H��v�k �+��v�̻�X�G�|}�(��{w��ju=��5�`^�ι�Sɜ��]�8��uNߚi��]3oA�8��x�O���A�����M5�2X��!�a��p5����D�I/��+�Q �*� 3���2
M	���pq�ps��{�)�9?fM`��%e}�Gp�Z�jӓ.'$�Xms��_�%�����|>��[�}7ҭ���f;R.�I���2�˰�,�x֕�MA:2	���6MbH1�֩�d�1
�>�o��8h&*D^�8����?P���ճI�[����<����S�\t��u���l���N����j�Y�2H�l�A��c�u3�/ސ�έ!�q�$�2�E"��x::�L��(Q�@�_����J�(�GQ!�<_����Y�:p�E�&)����	%�CV]�1Au��4�A� 1��=4�<�x7���Y����I��cV�I��M=XیϬ�  S��X�z�#�i��`�9��8�@tl��"Gϊ
�M9rS��´��M�o�E�-+�f!�x�S�I2��U:E7e�1��2sR:$�1-^vtC��a�$I��pd�r#��b~&��߉��ʪ}@A�sl���*���̉��/F��6��<�%g���J� �0֯��b@ ��[�C,����/�����܄���iK|C �P�����1���`On����$���rLvV��g�D�;�F�#y�	�S��i@I;��x�3��d��|�o\�箙H	�K���JF��_���t+��Ol�Sl��ؑ���j�ɟVu�:[M_�?�W��nW%N���i����y%{9Dl���ϕ�R5���"�~����q~�|�W�:_����������Z����4�Jx+����
��Ӏ���㌟�\�J�_�z7��fB�S���<��#"�-��y�0'�֕��7�Y+�:�w�j��B�'�R&�W�t�񭚋�Xm#4����f�%�V<#%3[k����
�f��P!�{��,R�����S���3�=%,B۳d�aY���21���ӽ�̒�^�Hp~~��(W5��qŢT����:��m�t����c�}棝#ѩ�x��Ս��н��J�"k��Q|���Y�f�z���$����#H�i��B#�A2�A��QmM��TR0�lLDs�}46�\ra����FwաT��(�b�$�EY:pPI����^C���n���V�K���A$|��#��A��O�EkD|[ג[E�jI�=t�LG{�ӹ�O/M�ƀHO�м��V�i��8`��w��^AF{��<�����r}�@)���!r��D���7���ퟤ/�+Qrr�y8c:l������~�g����J.��.hk�H݋v �FQ��G$�[\�[��{� ���a�"�z5�Pl2_��*�C�G)��<U>R)�v�)����U-�;1r��w ̿gK꫿
~Mh��s@*Yvy(r��H��b�ƀ�ʜG��������+pr�I�=��Չ�I��bѰ�V�8�5�y��2߶�tH:�J�<4��r���5%"]���+�D�Jb� "��`�_�a����"���>�*��nx�tRa��]� �ab���,z(��N��[�6+rc2��C�0E}o�����@�e4sJFb���<��u���t��D��hO�7)wC�+v�v	krǸ�E{��[�S�y�W�o��$���:��m����5A~<N{!����"�촹K<j,�r�]�HK�TNX��`b��%g���k�� ����@r �I�^ؼ�ƻC���+����7�ޚ�T�!>��)3�yt��cLC���J1��%�X�fr�t!��2��ϊ��bf����~�IC��C3��P��}���	���N�σ+%��6�
[�2���#0��:8!�sgH�d�Ys�LS4��A�諚"��Q%�"�p��A���!����%T����keY_��=2��g���Ħ�x�Q��Ŝ�
���d9�M���v<���
��B�ERIM;\��h41r�8�^�sA��EA����'l���i�<kD[Ѵ���7�P� jV#\p�ǟ����|qM^�J��.$R��U�g�.a$�_oX���s��jT� ��� �28�o�&�Ob�L$�ɩ]���xS��΂̄�dL��҄v��w
Ņ�H.�[VidQt��0~�ۈ0�a�%f��<����t�:��^d�x��4�:nR���7ɀ��3䧍�-��~T�H�̖�u'�+%	�\�c�p�Ȉ�Sk�i���c����X�aX��q���bǫ��@�?܁�U>��Xu�[�e(����yK�2'�0�`���@=��� ��V���S#�-��H�x��Q8 `&Q�U��N��:�:�]�ⱫE*�7�낚�E�X�5ԟ�l�W$N�iÈղ{�ce�@<��8X�c+2�Po�X��J�
.�'4�[{��K�i�vK�`�;}h��NH�MB�y�9ᒭ�^��y�2W�#?Ǐ����@�ݤ&4벶x�A&]l������Yۍ^$f1+X�/�����mf#��7ιR��0Ι'B%[	���9�1�<mQd_V �*���#U�j�7w�e�xpAܔf�Ħ��L��;��7�@E�{��TPԒ1��G�.������@v��������+=.�0��S�CÓ�t��=�m?S�p��	�m>I2���f��E���fW��X*�:�VH%��Mc#�xj>��1<3@(�tP��c�Z)a��Z�-I�Wt)�*�F�}T;)2�ģG��{���㌙va�=bhYy�q����U�qm�9@�s�<�z^j�5�>2ٹ�X���ҿ�Z�s�o���ڻ�>����gnL]�L$���ژz���>yj��/4rC�,s�� �R]�K�K`~ .�����r�����Ү�T�}���5MK3�Ij#��t#rKDI��;�LU	�R�9����n��'wx�R���,x�Ƕ��Ljf:R>lz��7����5ݑV@q�s����&;�8��?��?ZK����%�aA[�Y��N�����	���m �U�&�"��8��֊	�ms�'Aq@�G��I�h��12n�s��.�;�"��֒`�H��	jn�;�=J�~>��g;H:�X2��9nc�fň�	��]����v�o�6A15s�l��<C���><gb���59U�ڳ���)�w��5�
��-�T"7%pw�)���P�u4G�H��&L���Dv3ɑ�B~���n�������l#�X�8�b�3os@J�l\
�UAa�eF����Р�:Ν�qR��A�x��4nqa���FH3��x\2�6��-����H�ԂYHى����T��M�1�0'x�޿K�����b�(-p1)���5�G�Ire�]&�����9����U�ʃp��04�s�+�=����1������NwyQ��yNX�E��#��Z�ZHd��WF%f
u��b��H���?P���M�<nI)��7j���g�7s���"{��D������˨�{���L���������m]�/���,�Hw�ʜ�&�wR�G,�8̓�&Rf�(��EYʰ���F�\� bZ-�m�s�R�B�A.�8'���&��g�����(�o������䰡X�"5�,~d��}�S����2f�i�*	�,;h�5)af
%�~;P�^��wmE��18�n+���u|>��x�F�U�;���� ����pz^	8��8<e�\,K���1p��v,�~��3֖�
A�$U~$�0��!��a~tX�oj|���9o�^�䍭�d�u�U��v�0VzT�ZP�D�KG�n�E~���f_��İ�
�;iS�kndE}����uO�K��pYT�K��]���f�Y#��[B�ĳd��%��s�`S0#|��&�Y��C���(đŢ4�Oձ�2�_�2}�S�u�Kz*�V�ɵT�T�@\���xB��]8����?����/�/K�� �l��X�G�}x=�+�@/.Nc�g�!�j�����9N��@��֩��n�˙3UC�bOo�J5k�ez��]�|r$��x�:���R���Y
YC5���V����`�˹��&:�ᖠB�~�E3����5(����=*�S#�y����Z�Ar��<�O
F��� @ҩk�;|�Eu�ؖ��]b|n:"i��?δ5ǿ�bzR/��A����=��	�|�R?q���3�^v���-����ul�f �p�`�P��eh�L@U=�+K�{�ƍg���ZnpP�:+��{e��,�����r�]�.�w�u�D��<�Xv�&�^��s�J�#��4��t�ۆ��
���`�L�d��=�p�0��[�F"��|�&(�b�G��MP@e��2�g<��!��M��I�⪠�>�
���Entv+6�Y���~�P+��	 ��3�#�Ђ�z�k�ջ��u���Ak�0�`'���l�Ae����^^�ѱ1o#���'%��!hAl�5.M��LBk� ɻd��z��oՕ��D���!��/PfL^���y�9�}�魹=�co�
�`�Z,�a%�:�5�Z_n��Mwx��� ���c��riǮ�k,ҵ)52a/��1��qn`ߔ��w-���-Y����P�n8�dw�rg�eXU��/�|���K=�� ����6����ݣ歂sy�$�^2�ij� �'�a2�
�
��}�*G��a�������=�>��{�$��|�����0s��Mn��6��1C�rH��ąJC{����#^W��V���}���7�_5�Ue�����3��J�:���V\n������界�Q�h7~�p�q�p�W�9?�.��0[@ˆ��|t5���SsP�����I��]~��a%E�������Fj纋��Ty�����V��Ow3�FFFt��<��2�K ������n��!��e�%�3
���6XmE�����<6�Qd��چ�=�LpC<���wx�l����ع�]�e`q��|ih����B��>�S*���3KY�����f�&��FcS
/��@�˨7G��
�z�9D3hO�r�'�l��}�d<�>���k���/��A�����:�*rb����b��]�*��t���Y�K�N�Fcؼ��kB1����=0R��VH.S6P+�

����]	A�/ydu"YQ��ͪFB!��� �"����nJL#�"�Rk4�{X_�� �"�@ݟQ����f�Ko)8 �
td8��x�Æ�ך~[p�������u����B/���t^���
]k�Y ��m���l���Y2s��>�:y6���riC�l��A4X�j���ɅJM�Q�(qr�O���3�9qw����c*�ꍉb	{m���o��:�ޭ������8H7J&�>D\DL�VE�pj��7P��Ѷ�H�[|O�gۂ�O+�"��$���� �3㨵�`YCa�8�n�r�!��6������@^AS6PI����Y�T���3�'?8I̟S�x�� ll��>gXx�����%�hwJ"�f��
���}w�-怩;w �}�'�����f�t���-��c��O�2��7:���%��3�DW�1F�ٸ���0��3i'�ǽ������+'U���N�C�Wo�	�U�G��4���% Y�<�����7'�tx#��>�^$u���x��u�[Bӭ���Fe��>�]��0~-����ƞ�j�W�-�P�|������13��J�x�,��6G_}�����!�=����Dǣ��<�VU=�,�wЛvO�X��2t�9���iu�T����m�I��`'��su�m�A~q���s�������Ƀ�#?�7%Pm��>�X�gۧ���9�O;��?���
�Ǆ�y��o5���F�wV*�7�P�5qE)���I��E��� ����di�=�S��%�j�@�ƀXp>�7��Y�siD	��i$fn��0z_�Gk����ls�O��v`h������	J>�ҩ����!��V
�h�"�lb'=�pZ�0�h]� Aɳ�p�-9x���,+B�UP�ڗ鑀�R>�գ��(�L�7O�9j��K�N/;�ܘI<�I��\��x5��<};�)��0s�&��:��Gf�z��iH�
�-m�K֭��zo)ǧ�@h�0��u�'��
�s7�ApvrE�12�M��vR�A�2լY�*u��1��B2�f�8��<E�dp��� �?�#7���P?>���wI�ކF݇j:���7$�F�>TM�=�B� ��F���n/Aʖ�T/R1�!⎡�˦����%�4*2w�- ��A�w�k�f��k�� ���� o��9�h���R�a4婐k�Q�:�+�y.C�P|QVt`�8������]4��1"H�i3*Dc<����?}��_I������ɛ�:h:u������G��Bo%{��/r��������i�N�
-�|*��	������*����Gd8.&Ő������l����(�.���~@�%���[���Yܪ�6W�<��n�����TJ����9�/�5�I+�xA' ,~�������M�RcVTt�A�x��u�?�&u�ȿgNx!8;�"ű��_5�Dg�
 �,����b~l��!Ƚ�2��y�ټw<%��
�=ݮ*��@����I�Aqiw��S��tN����M*�6ޱq3j����?���R��E6΁�6�=�H�kV~�:��=�Es��7g���" R��3Bɇ��h�~�3i�RLB�/�e��I����|��ti٩��ɛ�.f�;B��:Y���8Н�"�:W��»q8�+�D���
��2۱6l�W����^�p�m�Y���4ɩ����I8��[��4��&�d8֠�>d� ��M��s#�.���ܤ�=U,��tes�8�]�C:�_4����n �n�ˡ�<T���c��}����	NG�pa��h�.�o7�92�,�"ѕ��N�Ϲ�}�m��S<�j��<���{���*��C��H(F1�]��:@�`���}� ~���3�H����<��&�޳.ғ�0��ѵ�c����	�eŷ<W���3(&-@��gϢ�Zl%�5Z�}����X�?�S�C�e� ����x+Q�\�f>����	��\� _��X2��WCdZ����s�,���q�C�=`��upV����&�NW^y5���6nt���;�M�J|C�-7dy}����A�>�mIFìڥ��0����Z��lS<��
�"�q���o�S�i�k#�gЛ��E��I�È��D�'�����%F0��?���6�y�|��� nU4�=N��?Y��T��8y.�wq�ωVkը��%) �a����NNB�ф�~��2:��Kx�n��q�?�}N��>�uw�� $=�!���y�wăYu�"�`(+ԁ�Q:[鷶��4�Lw̅���x��6G�I�ã�`'�o�,��RS��T�m{�F��g��8�&ᮩ��=:�����M��v��?Nh�j��uݜ��|
�����r�? tZH�l�()��ky�1,k���%I0�*�lC���4�ʜ�D�ed�\9�0��+�7����M�N�!�C~��!-}>�i���"�Z�~B�G��"/8x��v�a�ь=�	k�Ji�M'�*��z};7��O͡�Mi>]����w��F����>��͘q��Xre�c:�8B� Q�$�d[3���G d���I̪�b3
qpD+ٖ�"5gMHv�c䡛�G�-"�+��;+�1P �3�7'6h�$�HRx��&K�M@�Z��)�](�֩���l�,����O#&xkd����=�-�-GCw��=Zk3D�X�׶|ڇL ]�B�s��&I�H鮦/�'�$#l��!�A��t_nCm�Ʉ� �U�Q�EMe�*�s��6��h�}���;���Dn��a�;��q�O$�T�$G�;��[�ۏ���²�蕀��x7��i�dy��i��uh��*�r==pHߠ�Bw
�6z&��;��:��dXZ3�قj> ����O�J��z�3qT�A��zH�c�6­S�ߖ?�5��J���ۘQ"6�s�&�y�&oҊlh.pT��G�mTx��j�i/�'o�ͭ3��X+|�ڛ���O�cLsD��ba.$�����w�wj�˸[�)o
��x�A� },	�[I��7Ν�S�¥*9K��S@W/���`�f�j�h�Hх���2�ׅ
�Zi����K팎֑E��[�͇�k��2���Yּ��%E�6,�둯��,�C.H�Ƚǯk��}Q��Z���h|ȑ􌍱�H:���t5���5�(�
3S�Z��
(��P���#����ap�{;�P��0��b�74k _�-Iz�X{���Tl&j����Ǐ���K�ồ2QqL�:��y���� <�N�~<���i�VY2/^|��n[eu���K�j���J����߀t��W�b#-[\��׫�p[R0���j������1���۬��VZ��@��ΪN��`�P� �d�$�v��,Ad�X�/��ޫ}��E\33�>��
ȷ�xy�s��F�Ĵ�[�\8s�J�u����~n)���7��|"˵���A��YW��'�c�����{u�-Na9D��=�^9�DV��U 9���Y0��Ys���!/����59�ܭ�G�I��܃P9,���K�����^>#����oP~��%B,P�}�K�~єy@N��^���B�V���_*����s"-�b��m�Q����K#�z��Pᚠ�p�����^�v�[��d�V�Y@.��`�x�Zٔ%�V9��^�ao5a�C��N�MV �@��ģ����cT6��f��s�Ŝ9K(�r;JlOLkA;�v�^��p��pB��Q���Ϊv˂�]�0V4�'I�;U�qA���t'�gm��?V�b�o�\�"G1����	��r�@��Zz��'nZ�0W��pxմm&��ߊ_�G) ���_���b��e�{�OF��X��O�f�=jX�,�%�*�p/ф�{��Z��F���}���'_�� ����{�r��Q�|͟��!���jԶ,,�Ko���^��'��@��Eg���*ʻR[��h�Okf}�J��@�
X������?Hx�}|�.	��j�6K�"HGG�����B��I� n}��zt�&F���q%�;�$�q3�n@�k�]��q)��L�ln���	��I&i{b#�CDO�:`	��}���t߯��y[��