��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pd�Ύ���yya�[53㿅`�@�r���m��6��n�GW/w���Y��v��z�`����L�2'��ցy���3�{>��Ŋ)LQ �'��nX\
`xʈ=���q4��b�3�[ĭP���S�x�l�0_�>�:5��r뽳�8n8�^��}9헹|�K{�-���`��c�Ȅ�	~�q%O���A��� h�3y矰И���%;Hqj�_�+��꿾hz�dG�M��})=��nsB
�:�ZJ0�2B��4��޴�T)�o:���g�w|�N��H�''}=~&7W�؅yT5);|��e�(c|m��J��H�����vy���o�"m(�ޚN3^�ȕ�Ŧ��r%��'s��T?��,�b{�|�����N�H���:9\=�:�T-A��FZ��{��,O�/��S]b&XY:����S0�<m$I3ҟa�1��M>R��@�5űM�7�2���^���
���aa`�coyH4��t�,�X!�
W�J7,����Z_�ͪh�0R#� i|KY����	a�ߟ@��J����q�����<"����c�Q�f��¢��H������\玈��f_�[��7j�¨\3h��1@`�~�O@_<��/֡)�tLX,DZT侮)���,��(�҉kJt,a\�/A���>��׹���ؕ�vT���=����u�Q�H��9��5��=��+�,�w�����k�iİW4]&���pՏ�c�<7Ә!�G�mN��(���&Yښ���ӑPT_�.��,��T�V�������漀��eמ	�7����0��,��g��k�gT��TS�$�Sg�cTL���_���'������M%���by�JQ[�++�R�܂�mo�Maž9*d�H��S�:�*8:��mSn���U�I�_bZ+�ω���Q����D�^3`���uG��C���)vS���v���:��[�i)�#������T�3C�<��v��ܓ��}����V��~��l���cAdL���p�$��4��>)a=G�&�i�=)&�RFF����!��KιBb�PV�T����g�P�#'
��xUl��8�*�z��\��黿�,�����ߦ.'�����JӤ}�����#���<�*�hg��|kph����������a�k�m�fhˇu�z�2J��G�"gX1;y��:u� jE���]��W����c`|��K���Zx>�9�\�M�=�̡�P�FKWo����Qy�~Vq���`�e��D�`��q���NRg���a�o��! ~&Bߕ�T����7]�ɥM[�;UF�!3ǩ�I������f�
�]߁,��4������J�䮻�lׯ�Bx��+����>����Ξ�@�k�����G#f��N�SٟPz-f�y�����|?�A�K.��D4t����*�DT}��Ʀ�<L{�Y��n]`�簷�@��*q,K;��1�P�KӴ¢��k�"{�di�cۯ ���H�*	��b�,��6�B{�G�p�a�~��6����5U�ޣA��N��`Q��I�T�[R&"(j�!���� 5����զr|N��'##��\�|S�:9A�� D��j��U%��c'��'�ޚ�_3˜��T��wٳ�u���7A��7����;�45��_��m��d�%��(���q v���|S_:)��G�ρ����=�^���Bǡ�4���ll�Xj�s��;F�V�;�fn*{U����JK$~gu�S��l�qt韐pf1�Q���k���P���}���kҨ;0���x&@��O��ϙ�Â2@�\3�L���U��u��[��g��C~ǰ��E$起�,G�H�����SSF�Y=k����0P��_/0�d�߀�W*=��o�*� �x#���b����X�]���I1N�,�42J��7�ؚ{I5�^�sM�7$��4�-dr�u��Na��* #*41XX`Ҳ����	���t0�����bpn%ISNk��զ9�<��5>$@��6�������j��Uهy��Dw�>�3=���I#�|��h�Gv��p���e��j�&��bg(hC�Y����n
4���*Z0�V8Ѫ4p���%ecס����5��te�J���0B辖�-�Y���H�[�)�g���|��Rɟ�2�\�Eb�0{��?���m3�;�n2|n��0^�d��y��=*j�8�2;�4�T��R�����}4촧��7�o��.q�|��n,�y.�HCR��B"�Kz9�}lg�o#��T�����X���#���UY�E���(>�Ӟ�Cq�*R�_�f�4��sJ��2�u������Q/�r/�5�A[��C�-db�w��"X:W�?ukzpM��
p?[Y��:FDH-	̠�ĨI�4R��y��A} ��u�ֆp��nG`�ڜ�M���w�?^`�y"[$�K!E�ơ"���s�5W0E�FU(��C�[{�])��^"n`h��Z�	ŷ�0�Le�i�Պ�&~Q�bEw@Dk�x�=J�=�|�.��+�E憉���l������L�Ր
�<�[b�Շ���?+�Ol��0��VHHu����R��x@	�.2N ���J��kŽ�s^f�Q��sx���jS:���MtV�S��1��S� �
��\��8{s��:�7D�k�ed����WQ�]��1;�
�Md��0��X����哑�g�?$��#)�>v��=5� �Xn�g��������L��[Y���d��췬y�n����=2, A��bc�����,�o
�����D G� B��N�,&�0d���i��޸	F`qdR �/5�c�ӥ�Q�'.Cdѹ~�4��_�ܣ��>`>�f~^�5�_0�Q��݆󤳫�WE|f�ҿ��Cl,��țz�ra#�R���	�j�F���nK�%��M��	�A�H�q��T���d>_��Q� ����	���h�U���v���I&����ذ}6젶/���MG���K���|���A���3�l����e�����aW��}�6�ʊ8�]k`L��=�o ��/��*�j<GIϴ��3�ˍ��$je6��hi���m����g�;C�g��c��b�_ͺ]�X�{�=�*چv�sj�'�&�����X194��y��C16�����D8��iE�G6���/�hsM��)�) "��}�It�?���8LA[>3����Q���.m�lb�w"��w<`�k|8�[��ç �x�d�O}�NIm�4|��&c9mg�w��ʤe���6-^�PH|;��+19��_/zb&�߿���i0d:?G� �x�'��rn����X}�\��8�ߔ��,.��L������;Zo�O}17���:ؗ����A@-h������o�r̙��[Q�R��9�a% ��+�3A�� ���_+X<�*L7˶t�7q�I&�����#'�i��Yܸ����!ȇ�S�$�B/!�|^��{�*�V4@J��/��z��U�<��K�鎸pSj�$����\:V��MH�R�W����ekIR���U8) ��f����t��S�q�`��ADI��b����z '_�:���@����u�+Y6�Vu1 �u�nR{�?L�����Cp�{s�a���Z
���Ah8g��x{]�	|�"�h����|R�e!���P'�PJ����tF[�%<�j�J�(.2l|��;�Ҋ9�-�IK ��@bɹ��yҚ0M����D�8�f�'ҋz�o�ʉz|���[�"��Z^3I.d�jX�?��nSǥF��80m��d����j�����ϩ���c��
(��K����cLݩ�9!��ף�Xrr��M4Z!��mW��=�ʞ�����v3r��}��(���|=Db�����Su,���<�~UPO��.�;�F(����q�)ȷy�G'[zt��:�FL�����'�������A�f�@ �����ΥF����5���M�|��0ǫC!^R�����xw�Dz�7�|?sT�,�v��5Ĕʊ�fε���u��@�
�î�e!]&-�,��I`	TIR�)�%
kIS��L�ןQ�����T�ca���fv�([�����Oχ��N�
"gR�3߾g�WoU�åa�:�sY�&*�b�2����?�-N�J���ci�FL��fƖ���6Γ��� �����ȭP����Y�8=�V�ޘ��S�&S�QɄ;��z�ϟ �nF2��\B�����o�Yj�N���9O��_r/�
��+:�U~�cH��K���wӦ|��T���Z%f�]�2��_]���b���ˇM�[]�k�Q�}��7�od��#��y4'@c�߹	*4����'\ۢ���{��"��_�U~8�m�k6��*��J.M
�������L����M�x��1�K�=���T��,=�ڜ�����*��<M �kMP�~̰��Ӡ�Fy�\,���G��N�>\��dg\�D�����t�NIbRcp\Km}�T�I�b�'à��[�\�@a
���*�g�1���$��X�k��ѵ�H��7�Ge�/U§�@�����
2ȳl�0�N�~0l/��t7
Aw>1j�1Y��ݥɸ⃊V�rC����-��<��&?[����=��+��!*Ǔ��{�<N�w1G����� �~��ܜ/��u₂u�Z�5����+�6�Q��DH�t�W�>���f�p\n��̳���i��X���W����E'��nm�IW��W��f��Ρ<>�m�gM��u���cjޓ1}�Z��S|�i�#jM|������k�Jyk�_���bfD�7��-�Z)U1�|�<c�M�㤒�7fh_N�<t�eT�<XayG�;��E�M�QC"�xGfk<�?���՗*N�Dx5pd��_M���N���e}��	��6万��Uѻ:�1�6�����o�!�m�5�8\��p[�`����G!O��xM�*j������zZ��K�)��'.�%m�ג��2��D�ꯣ^V�C����?ф[BN�����%�y�8R�ĊD��OC�����<���5�Ihv'���B��i ?�� �u�����rN�#
��V��]��Hp�B��x�h
:�50\64ɾ��yĶ�Q��4�[��b�Üf���-v2S��������3��C���NO2KQ�Y�3�yN��|(o�SsM�1�M(��i�{o��Q\'���ƀ�2-�=��Y&���{;Y_er�>���$�ָ�y���^���F����.��&��&���>c�T]^����k׼�|�/�����oR3Uo| ���Nµ��ì�ThDáp�Rds��3�4&#t}pZ�`d->��1�8� \6�d�>Ŋg�<�ڴo��S��gb��}�}1	nJ�I6���T8bw�[��L���k>�������0೒���%Q�^�d�Mvn�����h3�������>8���!��!)�U�N�n���sw��2 P��:�pZܞ*Q��P}g��7�(�]b��h�7�}k��LD��k��)�����J��9a���H$��I?'ңm�b�D�>�J��ec�#<E/��9�m�5��*R�t�4s5E�m�n2���u2ܴ��ܖ�g�~6������1$�^LV&٨e�B�?�c; ���p�h��~�W�i���K�C�HM�|���^��!�#���|�S{�
���r�6�%�wնc�K튀1n�=;����R/w��[����.����o���W�T5���Q��Q����R�E���UC�Y���`��+��lc�{��:Ҩ>��=���3����ֲ����0n:b��U<���G�?���A����#R��r�C�������d9�����K�[�B�o��+
[3�ع�C���2���M{*���d�Xm�e���+��-F�Fj�/T����oչ�;�ɢ,qS�	�*�}YښE�h˰���Y~�������i�?ͷH@ȯ6�a��)�����)U	]�A��o��u�� X��l����Mr�_�u�b;TPo�n4��9l�l1���b����?BnO���ʳuy�P�s�A}v�xl�cRi�����
���D�}|B�Q�b� �>R���/$���~/��~ ��B�K�C.���'���h�����r���e*���~A-��#�
p�%�әn��~��T"O�.���p �k;&�D��B�;�J��s��/����(�M��ڡ�}��갥�A��v�fЧܾCJ �C���Mi 6����m/e-2�d~zH�:A�T�ņ��x��MŃ:��&���"��Qќ�<x���ym�cj���r�����Ex�A������w˯x7�XV�ѝ/3-�G\%u;)�-�U�0��N��Q���c�-�2��椢��A�6��0�hm�t�e�;�����	hh�����Kq�x�� r��H���[x�T�&���7�i��xf�����]3�Ң��?��O|>�7؍�z�!��t�΋䁙�t�a��'_!-ݟ���'��f>��p|��>b�����|�|#_�3�5�$o+
��g�L�����Bg�����Wzxх����\��'���g�O&���m;?���s�0Hԃ�j]�>^�� w��yB��ln���k��� ��o�);&�NI=�[d�n��
 �we���NO/�FQ|*zPy)��sFa��D���5����so���l���� ;�j�;5s_�1�2���z�;P�f2'����w��`dq���e)������+�U6�%����7�^���Dcf�>���%�z��@x��u�,�(dĭ�Z9��͞g���^�����P��DBw�Lb+ �5���>OK�ޡ_�(�9I�C
S�l)�3寏�O?%1����Cmo[�lYת���Ҋh��L"���	>bT���8�Zʊ��u����	�H8@�Y�~I��>���E�Ϟ}�dn���/�rJL�8Yc( �jM#Í�a8;D�����Q��v �x��wɯ�Y%)ւ��3����:�݊�_3	& ��m�Q��ҫ�ZI5E���hf��.�@�����3��T��	v=?�4�A��a4��Ī�0e��霨.	��'�7L�BM{х����� ����4����tM̕s�ߥe'�Z�%��'��ܻ���e�@���yB ������%D&�:�=�X�3�m��gg����%o��& &JH$qi��� ��Z�(��]٧2;uG���Xl06�5���?��/��
/�R�q��݌��$>�tOkA��e�n�{o�.P��|;i�N�Z?>J�s[	�z��ڹMO���|��0��_�w�//� 곞J�B8�$���Tz�/Ц�ᴕ4�H�Z�)x�	_N�2~��ow�Z��b�+�P	/��ɰ�cuFq��6�N�r��oh�T֬�
T?13
I����³4b]�o���a	�>~ͬ%��MkK��R��d�0�Y�������n�|	��66ț�N��axP*�S0!����Nn�ؙ�	m_��X���f|,����D߿B>�:���V/?�t������X���B��V��cs��Au%�7�ٿ�R�HE7�p@`�(�dD�/�)�pٕ�,.+��G��n�B1�w��Հ�F�)����"�14|�+��C�,?yzӵh�/�{�C+矩5{֣fQ�1D����xY�KF��3��\�""�/�D2J����d�G"4=��� �@Vo�Cv�4NC��S����@fY�k�2źW��U��^RB�������Y!-�>ղ"Y�T�R�����K��� � �
7��ef�4WŗHb��ދr�N=kE2���|6�eV�&Z�D��ܽ���S���f�Ihx �/ҵ̠۳�s���U�[���Y��7�v}�B�R9��Z�	�����&'B��$s��},�)�S��)��G��(�`�Db5�3��AU�@9>�tT2�ƚ�F��m}ḻӴ�kB�lṫ�J�L(fń}��=b���u�̥U�m���:�j@D�@?o�@�)�KT%lzOץN�a$2��GTx�$��I'K4��I�Tu�� ��=q�q���a�3l�],y�)��C�5$b��Uw�j�Ȭ�N�#��txx�1s�1}���eʂ�S�� W_5'o���Ӱ�b�<1;�`��R<̥��8���&������U  �o����$���}(s8J�}��z�!>�8h�I�(2U�D��l�j���N &v�4+�|:�g�wB<�)`/u��s)2W	h�I@T*ȋ��~�IڞŻ�ۈ��1/ꛯ�������|��q�4�M�P16��۱��Gj,?/4a�)��]�f��(�Z���3�*?��q�'Й/N$�_�?��a��/�����(��5d��[|8��E�Q>T�z)�;�R�<zw
8M��� �<-(A��5��]'��[yc?�X�M� ����=���Hf[گ:��x�+�<*�) ���z@Ol��I�0��K���N�����]`�$�}��X�!���N�rA�MHj�5�qj&�嫌o�A�0����}%�Z3�P�Y�e�c����"zE��QC&J#W
E5WQ��iI��X�ݿN��	�#�)������۰@�]����!�D�Ge�H�����Yw�F�� ����L<2�E��>�B���'�	��M�t�׺*N��Ҕد��B�l����3Z:�����|,�a���!%5��
J�w���oɄ94/n�cQ+Pq8	,��e����H�>f\�����2CfN�D��S��Z����w����k�X��W�17���l���D0�J�ly5;z7^�j�ڤ	��<5=� ,�"���a]$�����^���B�6�)t���f�s��ٛ�Y����q�� ��9��h�H��ڱ�H���B]�3�� ����TOhۑ��`���ǢɕQC���I�`��@t���;�k�[:�?
�����o&}y︠�p��T*#U����K��7D�-p���pO���
��MC���N_����>�̋�A����R#Du��>�Ǝ��,kV���qA>�^׊W&VOE��(��v��J����P���n�|f�oT-�9�3O؟��Âh��U��ҳ��GX�%p�X��L$!m������&��.m�^�ǚ���^����[���H�s�P̯�/>~�o�	S���= ���i:7h#xi������dA���~ӟvF�d��nz�h!��H݌�L��E&T��vI] ��WjX��
c��	�_��!K5
o{����/\�SQ����P}�k�f׼b����Y'����J���<�n���F��Ӷk��󈞕�g(��2ݰ����N����MW,���ɑ&�Q,gU�r�*wq�b�/
��Y�V��e	���m݁�E�ޓqg�a��E.,W<GDwh��K�I�Y��x���?~��3Y$��^�Z!r0��G���ݢ�y�3V��}�ݒ���9����#kI0�v{ϰ]� =si �\��d�_��H����%2^7����w^�V�;�#����!�ƨ���l7���ޞ�q)�aN����l_�4���j
���\9Xc<����.>N��;"T���)>{o��תw�Z�<U g�-�(%����h����,�d��W]����L],_[�:y0k1N�]��X/������%�I01��Qʊ\(�)�k����>_�u���� ��CaI��c�	�~s�����s�1�q��u�Y��F�?*I_�9��R�G��4_k��'�|,�e�!|b��0Y����Z�_��_U�G��GN�L�NX��mW�voA ��E�������>D�*�-��/��d5
������"����F��#{����%z��ޥ˝�qB�y���'� h�x�vn�+������eu�C�"C��(�?v1|-U
��R�d^*y8-�w4�O�E���g%��E�š��DrA��o�/��u2�o.F�=�6�|U�;W���7)YȢ�E�X��-��W_Z�A7�x�c���N���~��Anq��
� ���-��8�,x�t<��a�1I"�}X:!�J0|ˮJ�d�}�,G�X�OBB��	����v��G~C�����u,�X��B��EJǽ��*4�����¨*�V�w��@T@P5
<��x��+vсA�*���_c('Ԋ�Iq'Yl>����@�|�1����۪�i����
�����t�h���%�|;�șS��x�h����%s3���zl�FU�BБ�0* ��#�����Yi1��EA��x2��aE+�f~o<������6��W��Ti�AZU�F�'�:G�=����Ĳ�L�]E`����
�퐰��:o�.�}��al�G�yE*O�����f�}�ہ��:�l� �{JUۙ�o�l����:���^?�ꓶ���z G:c���m����A�/���v��_[���w�ˏ9~dF��N�S��#��%r�c��Z��X�1�#X�Ԍ��7�_��H���P��wr߅�y�E��0P^�*��qW\W�f��S���D:��{>�-�9K��sH�ǔm�q��-�L�N����1:y�B��'S�ٮ�e&R���>��������o��&����b�W	3��7aX"��J~��We	Q������� �����w��j�'��-�D2��'O��,�L�ϖ��t�AĿ"����j����^��^�����Y.�/�%��%���25���R��(��s0LQ6��}�j�x�����y	6�g}MJ�˭���P
����V�!ε^�?�B��:A%g�]D�����6�^�@��#�ԉ�׾Y~��n���-ڼU� ֛B;�f9���Ɛ���q���;d3���׬6x%i�Nׄ���uc�1��w�%8�A��uf'7g_����'A�x �g���_��u:!!�#[�	�Gt�岭y���@3Mq�0��9�3{ޅ�N�IoF�I�UY:�/�R��V�zɣr�����Vn,�u{4K�m9+#w��<��B7���f�	�}� ���}�������� H��P���t��㔡��^]_rxI�	A����Ix ���W�a�L+*o�e�� �Q�k����`��$�o^�b�����]X,��$���E~9�U����o=�R ���9=c�����L��u|���^C���T@��st3dsX7\v��� �g^T��(�N��]��hc�r�����-�M @�W.����1ٛu� K3�b�y@$����؏ �)��\ț�Ya�[��Zȿ�2�kw���6�)V~���d�*(?���u 