��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&Ű��=�b��vT6�4��fWg)l]��@��7�B݂Dۉ�{��m"�hIΞ��`�$p�}z�Ҳb�ZV͕�e4�NU#�%���o���j�!<�P��Ss+�Z�rbN$&�a��A��4��zJ¥��	�����5Ӆ��ar_�ЛiA��,\�FY�et���'��W~��b(���u����Hg�Ζ��M�����h�ڃ���^DY�v\X8Gv�j�&����<��^L���c�|��AY�~e�R���k!1,p�R�������@2T�!0�(Q^���Hwe>���k1U�,���{+��~a�U�#~~��5z��%u9�N1�3�ZZnT�-�*�!�n���ؖZA!lV�#���q��H�
���{��^P��1�|T�Ѷ�S3l�IY�N�[f~"��9�ѻ8هƢe
1i >��R�����h6%�����1�v��s�e�8J\����O�>��^�Z	����&����aN�{xU��*��F�����8�}��p=�����Z�"�v�-/�P.L�����d�G���Z�@�Ё��E���5�ô{��5v+u���s�+�/C��o ��\��K5�t���D�'�RL��Z��U]gh&� h��ʷe���y��JjA��X���b�6'x����b
= #j���d�1,26HG:�	z��K�Cd$��LJ!@�P'���Lw���ӗ�@r�b��&�&Y��2a�-8K��t�<0�8P̮-;^�ot�W��K��7������ڷ7�_��2CG�!�`8O�I�S��	
�b�ы�Fm���Rr���t�/k�<��ѝ�]"��|_[PC�\��VG�a�@�JR�����Q�q��@���J!��]=^FI�00���~��,�ڑ�7f��ks��ݨY��cbm�ƫ�ң�,�����d�e�Zh>�F�ik5,�����!�������ᓛ�u=4kr	�����zL��23)}M�9c!�D��-���f {o�gh���j�P�o=mv��M����Bei�R��E4	�}Ǜ�����[�SyQ�p��~�m\��*��_�Z=�,d/k������~n�4�i�����7�f�,$���5���W�+f�1ȏ����q#
�@���G��������jY���Ac>��E�=��I|P��x6Hw�WL�#�
����s�:�Z�DlB�'��޹/��J���
$W��C�b��]�<t�Jܷ/Qg��b��Es[b�/;�u���I�bGγ�iɳ�ZImܧw[�'9x�'�--����~���3
S��a���
�ٔ⪖`W�DVz<:�Xz/#zj����nC��E�ʠ�Ϯ�f5e��ь<�Y@E�����| �
�cE]��R)�/�����`��,Q�R��^���ab�
M�=6\�P��C��Q�'�[����4L�����p�4���zT%��Ӛ�{���Р�u����B�
�6*��,t C$����U{�A*J�9���yi��Vw�%��2νFQ��h�p>���q(c�VW�C ����(,(p c�6	k|NzȮ^��T��dF�_d���ѥ
�NقN(QN.�2*D�.|Ҁǔ���W�_3���?��w��O�ឯB��Ӭ���N9���!/\aQ��8���z��Z2U��r��3;�`;��0�w�9�:��ܺD��_���j������.�����ѷ�E��x���6e����O��V�ɻ�Kg:@/kQ|(����׍����St�>��Y����`�0wT{p1�����[�Ǜ!�pv1�s���ݖ,CE�,
��LY
֖"o.5}5Ov��;׽�,�e͗��7�[��Úv���A�t�_G��yh�n��-y�
-j1��jrܨ��]#��	�r\'/��Q�{T����q��`z�b�N����W08iK���+:%�xv��S�V��~�e&�Q����� +H�{�S7/Oj�\��A��Vz���~V�k;���{�uȯ�)�Ȣ����1y���P�E�d�����:�u A �7JS�,��O�}d�
��Y���K�ǔ�o;yr����Z�7�k�4V�ݱ$��G�R֧!� �>���9�#������E�W��[n*)���c�0'ǣ��+?�aYu�8�bw��h2S�fSH�3����m�X%A�Af�|�J�n�cb��U�~
��j�R��Ϭx$Ēy��І���Y��w]�����j͏� �z߽�X��&����LҭA���c>��W��J��IsQŃ�^\�9�v}-l�$.G�<�ْ{���_��.	 !o/�lO����n��E�ȁ��!˰ }�bN��f�Mk��=Og��� �>�s!��E6��GBaAB[���4��a��QRN�4?b����?�L�L���t����ҿH qo�FSdh�^?P)�+U�x`al#�Fʖi���*Oޔ3i�,��OT���H8��CH*��pΊr�Vl����L�O]��Vc��E����T����\|�����=
��@�~|x�׽F�ܗ��ht�k�/ᒢ�@=0�H�s/ 	�ᦘ�̫a���K��}	6l_}��V0�7Β�y�����>���,�|�dϬ-��I��Vȡ��V��[�'>N���½��G���X�зi�	FD�W�R��̙V���]|:ס�Z���N�3�I+�IG�.,���Ǘ5�]��i�v��QΣ���k#���1�tq�t�K��Z��jו`d�FR?�O��mݫP$X'އ��
{16�{3�v�@!�c	�ǆ���T��#��DԜ���XL�)V��P�ԘζК�`?�f>qb��7�OV��q�HX� �r���ϵ���eG��R�VQ�A��x�z�]>�@5̭	�.��~_���bR���!�\l��
y��`G_=K��A<:O@ƗMn�H�xM<C����b�9����R]�:�~ �J�YN�{íݺ �]��{	�<E3��V����.[k\��������\���m]{�Ij�_ 6��}����d
E�K���t8V���а�r�ϸg��S� |��$t���.���[`��ݵ��|xk��W⺽���Rq��:��H���:j�~���9r�U-�|Y6숕���\�Wk�W(��X5��;��!t{�V��J"M�� �j��>�Ry~�W��<��H\�RWpȷC�vE� ��l?�3�b�r&v-֧hI���FV�� Ì���>8P�*���5�]o}0��D�mZ��T��;�i����E�Ϧx��s�*!
1��jc��L�ˇ�L%ډ�����-��;��]hn0LV��3N�*O�,232��_r^*W��\y����).�"QfAb�ISe�T�;pۥ�!��!3�0񌀚�u�39VM+���-��Y�Y}P�v��Y��V!9�s~\F;c�0�OK��J�y���ݥ��Pk�F<����Enƈc�hH���z2bWSF{>����s��Z��*0/x!�m����	�K����4�=��N�;6L;W�l롿zx#�Nj{�vڵ\k�5�$TZ��s�L�^c�&��q`�9Q�To^�&�U��!kv'����"S	�bD
u 'Ѧ<{-@����k��uZ����qGL��!B�e+$��=?3�Ǩ��s͊j9peK@�X�Ȓ})[�H�/�i���-e��M5����4T��N��T
4�Ηީ��ѴE��!��a�ڴj������u����M։�?
)K>���B<���]h�JY��S�{C��Ķ|���i����.� v)���!Y���f1��,���Ev�A><;ldM��]�L�AIٱ��~��Q�v�;�Oe�K�>D�)���}q>�^j�� yc(�t{X������Pp ����Ol���� �la��fO/܅`����r0��u�C<��Ϥ�ҖVG� M�&f��|P�A��Tg6�j��H�^���y���Q�!��M���%VYX�� '��-.��	���q�i�t�G� tU�\_�
�2��xLָ�7��󅱋��7$���7BӼ�9fƵ��\�Y8���bA����������Q0��de���r+��m�z�16VKu9/�c{����O���-8.�o�@���̆(�gh� Gd�V�{��!�Zp�Q�j��e�pr���uyh�d]�k�M�����QE�W^鞘=�:��!�U�j59�m���pc��8��e�����A�V�s%��b�2K��X��oi)���[�ez1!1�@������rR!���($�[A�lʦp����j�({I�8vV�}���t�*/��{�n-@�`�{ȩ%Bt3����ʃ$F#�|/u���o͠V������n��?P�v�NF�)����Be�āyZ:n���(��z��\B$�P��8n����<'�)���T�nϤ'��a�%�uf/����TT�k�ʉ��b7�z�l,��9GY��'܏@�-4�y<���_� ;����8~l9��SY��f����N^'��p���wl��k�,\u�JW��?\78�� �eh3�H3��/�!kDݝ����s1��V�,�@ԓ��*���>��W�����x��q/�8�Ӿ�5,	�9'*Z'����;��d��m�TɭJ�e�]�y�vb�R,����ǳ3�ccː��%{����垧�@�3Z�&t�U��+dV��D]���U�D�S��*�B�u�m���K���[������[\d�7��.�	ߝ�cY�61��V6F�B�Tib9�H�iTk�6ą�"BY_X Dl�
�'ovB��c��8���|}z�+��$m�[�D�<��4�$�G!Ǎ��6(8���PLDc��"n�7�!wƭ�Y	�
ufW��&3*�����^��Ί��J�X��3�<�4�`� �Y˽�YѪ�[�n�`�x���RX�ӛ��F[�|��,���o4�d#[JW�eEb1��~1��P��"�N�PV����hh�N�O?�@?%�0��!^�i ����TF�h����M�O�$#@.}%�9_������C��^=g�$���?K�P���'������U���1����͍���~b\.FC�����_Ԕp2�}�
�1g�	TZ�|%�����̐%��i+���O{
�J3�/�V����`
�Cd=����?fp��I�K�<�Fk�̗T<�B�dН�E�Po-5�~ώ<�2�4�I���آ�X������K��kZ�c��b�6byw�>J(+W\Kx/���J���F:��a*\/��=I�H�軤��vY��i*+�AbgAMgE�Q��E��	,��3j�_;c?�	vw�-w�C���g4��&�{q�°�'��?�f,��5�ȒHgKqB7�9Tk��R�P��2B�X�1�׬�Ĕ�78lzH_JN�3��C�0���Po���l3���*�q5�A�kiSH���s���*��䏘�խCW�T���)�p�����#��N�����sor9+ݢ����i&sjfQ2&�`�tZ|�_ɔ}��ԑd�>���m
,�J>yN_�f� ������ H5{��1(���$>؂_����g�lUE�w<%�D'.�.x6���D�CS,�����[ɋ�o0b=���d�kdb.>��d�틼F�M{]��|��_e���z�ߗ�x�6Q\��L��Ey����G�Y��$�o��B������+�h�\策�Ħ���c3�f[�#���X�$'����S�T��{��?z�ޝ$�~ي^�p��N�3WF�M�H�eP�
���REC}�/�5�x���_���n.�G;��i�'���	-��|��8'���~��{�ܒv'�x���f6�EX���I5,Na�Y��$�K�L䈛|���w�?1(��B�Hi�&X$������%n�UE6�D�G�
ۧ�f?,UvG�D3m��ë(��?О���N%H2�ߥ�b'�i�ϲY��F-<��aɰ�����4�KĩGd}&����$j	�}�҂:��*Я��Y���i��+GAm(�l����MF��#Zr�]E5H����h�]Z��,��jU�}�}a�u�x�8�p��sl�v�S��z�Ȏl_�8��JR��;T���Ml�%R��2�fp�ӡ��#�8���&[��6����wciC6�@î:�		"Ż�T
w3���Rx7pF}�u�,�
��m<X������ڥ�,)|�f�3	�|텖�Cg(f����fG��`��j�D`˘QgZ�p'KMr�����L��R/ ��S�Tu���7�����|�[�0����4:�Ut����SD=�"�+.c�S"��%�!���I��rA�t��lU
���BQJ�(�<s���غJuR�d�n��%�V&[����+����v�\ߐ_�Ɔ_�:P��4>��eW�I�:���p
>�p���ŉ�����G�pkTTZ�.����9�J�@�XM���&�d)ϥ�ҍ|�xo�����V�N8��Ö��\���c?E5t?�I.�K�"q����s��4۱&8�ʗ��r��p���*���ġ[ɝ��7e<�����*�D<�0�?��2�ﰘGfk��.��Gp�ֵG)�:M� �����e�a���+V��H"�e�6�0 k�l\�Kwq8?r���5Ջ�^,6QL=⏔�7//���Wo�K�:r,�Hn:췲}��CA<d#ڜƠ�y��]^>��P��(B0[���"NVx��KP9��F�`)ǥ�9T)G�n\�Z=��6u�
 ��l�f��G�쐉=�A4��ene|�<ݥZ^_��԰@���I���DF��������x���nA1zVr?o.R���#H3��i���N#	�KZf�����U�u��L��m�S䶝���s��d��Hq�%q�����C�n�=��O���'ةP����hXk���-�7R4���]�Q�b"8pW�e�_�2����_fr��CO5���-��w�8YD���3k��4��g#��ÿ�.�a�ṏ��1�]m��BΑz���)�i1'Ӿ�S<#0=���{�5�L~�9lMT�75�����5�̐x]d��V���=?p����j�������y�̣D^�Hظ�|	�_��3?dA�Ʈ8d����%��NldD��3����ɋ�T�����]Mޒ~6=�,�)&w[Em>�{����=߻=/
�p����5z6&�2����g{���٠O@�.�̍��g��G��"��$bIg����D.P�H��Az���/`�ܵ�@��t����
�ٟ�6����\v�e�C�_&0�Y�rB� �����<��hk�l��
;����Q�J�~&�%�l��"�r��^C��ALc�D~��߀�2$�L�wv|���p��� �����s����O���ZI�F��͊��ɿqW�%Z�H���iw2���}G��9�I��P֣��7�k�b��e3-����NS�2��1zC�~>�-pY�ܜ�L��o�'�ӻ�����%�H}�0��pc??����I�"~-8���&��Bc��^�x�.�wW��,�^�s�o�>���&��� �=���+ =��%?����1N��o�\ �~[aN�-��86���
 �ѡ���.ٲ��6�;�&/aM��^�+�b�����%��w��Ś�%�vXD����(�|I�y�@�,TǪ|��j�6H�!��d@���Ԁ]%��<{=oH�?\�_%�샥�2��=Gy�b��O�祋���V��1�o�ξ,�2!um��
݂�v���WG���-<!��6�-O3����ѶUn&��UӠ\j�h���2��!=<��Z}[�E[��b#i�4�4�-��&�j�B,�w�C����h3"Ù���� \�X\ҿ�*y9	U'�� 4K�Rc@%gr�D��1y5���U�kʭLe�**�ϙKoU%�h2�Z�T,���{���_i�ݗ�b���V����E�
v+.�m�͓Z�������5�
#�����X3I���.�|Y����S���gZ�	 �A�2i�����1#r���'��RM5x]t�T�#���ES�:��Y�9_��N��:�{sWh��lE7I�׷A�C��ڵ�x=�O��+�۳� �k��M	�b
��xL���З��"��&#w3Kn���w����I}���AfOFu1��E���[�.5VTd抖�d<p/��&,�WȔ{|�ǯ�F]|��GjE��Z�OQ�pׂ���I�8H����'�7���M_��x��\��C��7�S�y���ۅ]_��������Gu�0�?�@���| �y
n哲�v�Q����}C����א�j�<��#��g�6/�շ�O��`J⍈��j�$�c-���Cgq����H8�o�e��}ڹq���Q�q$�į�h%��3��)eyB�z;X�z�n&���{M57�ܒ�ūC�H��l[Y�"�kh��CtB���-bF@'�d��16�""Yv�\�Q��s��:�L��N��}a���Kg;�"z�Q%�k��<�����v�W��N�ķȇN�n���UM�U�F�Z�eh���pR�ʛ�J��÷�(y�8��dϔ��8��4�hx<�>k��#Q�j�yQ8�;����xy'v�C����U,��h^��������u����2���4�Lٶ���uM͞g�_M逑j "{vD�ꑲ
q�i�yL�rˢ���U)7�lS�$�1��Љ�ey��B�w��p���팮^����>�E��A���ә�X�N�ŭ���];>ܡ��4[�-O�k��&P��! �q+J����L�qC�t����w��}˯����̪^�l�G��
|=Q���Ë�A���>"ߩ�L%�Ӭ��j��l�،���Va/!Ni�I�H)
�SH�E4q�F)��#��V@�Qs�����Z�w��>���8�^��� ����<M�moЮ�	ZP�b]�M�7����2ij�� �t�vpb�J��09?�#hH!R�_��y�SЊ��n�s�X7at�e�,��E�[%N8-�qHເٶ���D�r����u��;ћ?P���L�t�"�	� A�'\F��х��F�W��K��e�,�)O�fc�NFgJ��#Bg���ɑ�6�6�a���tt�x(���:�4ѹ@^x=�ڞgT׿�f(�YL~�hIR��b!Ag���f�*AYYV �
	^��K�� s�(��y�o0ò�WNv��_�30z<t�:�kڌ{�l�d�*����3�52���rS Q��o�i�P��	��� �,�_����%��(��~s]h�S��(�3�հzpz�5%�Y�[;�lt�]9��b��X|�hg��ێ?��.?~%�1�k\D$���.K%y���kB���R�I���Vx�[��ˡ�i���r��������1����^���[Bt��,F�?tz�_�X~�r��E|ٱ���1�'�!�,���S�@�32^Hce3S�����4'� ���Z`��,�qdM앩�a���b9��P�l�)V%�C�^�������뇸�pF��s��b3��!�ڬ$��/3�o�Z,c)�"�f`�@�Hge����X�,�p��J�t����)\�[<��{���J��(��)��%��p^��aMg�2�~��XwI����S����K�3-���q 	���
qh-�3�ԖU���:p\jb��������G�(�ҹA���4���\�c��J_WWLڑG��6���d���1g����N��8��!{�x������C����d����m����)Nș+��kG��-�Q��q��s���fd}�kEG} �7r_$���2��&�y���XX�;��B�:�� �m[�F�4�F�_����\��f���M�}i;�/�;��j+���\�G��{g��~,b����Sƌ�Q����Cq�	�9̓H2ˋ6o�.�QV��͹@��x��f���ȃ})�;�`z�������Ī9n�fbFG���93\��b���[1�x���^V;��*k�cd*?�^�i����4 �z4>��}�����\�8H}��,=�2{?w�fw���\O����vd�	����c'��P�_�>�#�AB�mHG{p����z~�y���H��c`��L!k4�x���]*��b}
N���fa<��O�+yo:��&c�#��	M�t�����+K��P��r��J�A��&PX���g�\�M:8�j��V_����zX�b�(��Yg7VGeW�@T%i��:Qy�z���P0Y�� ��7
<�����j#]jf� z;$)��\X��23ꡕݲ*�&�x��xD�� �\^Ң�f��- ~L1�S�(41?��� !�͍��dt3���8p�+5#x6LP�k"5�kq����z|j�o��9���D��xDv�2�)OKDh�g!"�Q8�V�J�`����K��h[���;_�ޅ��;xw��0��l�`q�lb��P�tp��S2m]=�-1���a[ҧ�p}#B�
����(p`Nc� &�Ǣo��Py��H�5)����m/QQ̥�]˩_>��u�.�u
�J�����9��&+�d�H�7L���2GP�ETM���/�6@�Sb��ð�D�K���i��E�oʅ�i�Œ��i�{��}���wG@���J��u�!��s!De�*�׻�a?e�s�|-˿���eDje���#d��EرLH^�%,S�:�>Q�~Z�(��%�,�~��u�E�D3Ө�M�p�TBc�\D��4@��O6�,L���r���5(���A&'��1O��\q�l_`�������$E���EM�]t%?�Ko�a͸Db���u�Lgr�`1���st�U�=��.	����/3�l�q�T�	��~��.5<��r�K9Ls��VmX�������d?�*q)��<�[u�e�)�g��߇���6�˟[��j�͓� ��@��J��7l� ��Ӯ���M���T=z��
Zż�[{ԣ�>S�p���&5��D�������
����^:BE7��ᯚo���h�4���Y-MR6;tQ���Qx�oKDb�����v�/e(2�Uڪ��O� ��#����D#�)ɩ�˝����`P:��/�@����öPaz����M*�U���$�]��U8 Q���\ڔx��Akf�<��ڠ{Ql��Q��󚆓~1������Dj��І���o]'���܉Hcv2Tc����% ��+�(���;b�4�����1��)Ā���c��^�Sq78�_�H���)I C�q)�~�{�J��yf���	
[]-h`�������J_y��U�n�)��P��K�s�v|W�t3������.��c�	��_z��U�R�����2��Ӝ�C{+EnX.�'ǽ�Cd��X�F���D!�E����b_���5!;��$�"��2�J n��=��"�Q�P�[]f��D�M�j ݗ�6�x ~
w?�W�
u#�Jm6�2�� �,�e@]�/Ճ�0�Ȫ�W��B����>����yH�1�,u%����-��G���5��-�j��k3FjNV@*.�KS��I�1-UBV�M�q\ﳬ�<B`�ِ�Ȟ�ɼ�;�W�u���s��f��Q��h�g�Kp��'���͝F�XUP�N�O[�?��s ���qw�G���ã��?T�vo*F�1�Ikb�pп��K��̀��%��3��F�	�8m�<���%�0�q�J�����~�
E'v"U*Ẃ��R���e�X����y�nm�g!��xi;0:ãe�2�l^�)D�-�Il?�~i�2���P��L�c|Ҵ5�]I�SE@���oBrT&�/�����J�la������J�j!y[h�A�p�巧#�����?�E������f�$4�y�	U�[�V2��:�wE�PȍK�\�A���c����d��{C�i��-{,Ps�3�{9�f�l�w�4���W5q���V@z0]�*��z�N�����]h6W;��j���H2��EtYF��J�s��c�~o��=��{��1?�-�G��)ͩp#;g���j�c��Y�[f�8�]ԕ�P}�)T��6y��F��Yu�EU�M�cT]B�(\ �6:G�>��N2��|_j�W���fױJRǐN�
:e�3��#o�9��	������B!�PCg�~i&�Kz�Z
J���߼Vd[�v���" ��eK: Ed��v�3�j�c؄��cP��"6v� aIj 5�88b�U$/Zr��x�pt�I�%��y4}����X-S�y鍵�"��3��j��J��zm� �vɵ���q�XF��T��vdVδ�=l����A5�F�}rt~;Z�~����ey��J�m��}BgF$�����X6�So����rF�V5SW�����B
d೏����S)�JEn?�Y'k��R0DS�|^��zn�g)��i�ؐ�"PJ1"�uM����$�"Gt�<qy�x���;\i�����7�;��8~_N�I3 ^C�"�Y?�	��2�Z���г����XsȯKA�����X�G"p��e��qq���7}�	y;��an�WSz�Rr8^R�+D��R?��"����D�R���=�!J��Փ�ߐ�J'f�${=#�\�:7���w%��*��Ǔ�~r���*A��Z�\,RV'x0��u��6����ŀ.���O��'O	k.%�:���[�/QE���o**z��u�YCI.̈c����wS;Iz�ơ&��Rq1+�XT��KC�d��7ڛO,����'\���)�=�����Q�� ��:ƭ��g�^�E��:��z6�j�̸���ş�_I�H��xnT��wJb���k���z�!�S������S�x�UxL�p����Zg۝��"�}6���^U�]��ɹf��qg-9��%1��T9?g5@ X�1:�=R#o�������'��GC��\*iy�o#-2��P^dt!-�gt�Z?9Z_�<����.%v�hׁ�x��.�쨼>0l�����A�;&��[�ډrĺ�S�8�����&���x��T���.��h�{"��h�ۦ����tiC���� ���z�y.O$�J����{�:;]����-�v:p2�B�n��+�`٪��{��K�&�+=�0� �|,����ϦǆREi��~��6%����F��"���}?�}�;$���Q	��u8�@lCs��oy�6QR�G@->�/����^��h�"��ⱗ{���9�:@{ÇT�Z��$�߀�(���`��AU�ܚa�r�$a��"�aZ��6wo����k^C�YI�SlyM�P�,z�Rp#��e�����������N��LQk�~�Mſu�)Rx�¨�D/P�m�#�1!��0��hg�3���<-��w��ԧ�""	�"*g��˹·�g��  �;'0�I�~�H�}VE%̓^��n+�b1D�&5�%MV����ǌ�u�ꋍ��M�$]�Ɣ=��g�����f�M�q���(��Q��-f4�����;�c�f�(;�]���^T9����X�p��\��0�c.��
q�+����q$J̳r�{�)38"���'Z;Y�S%���-��$��z�Xa���ʸ�E�yv��f�_J4���*x^��$��C ߈A٤��$q#��/�o)�D炽�_�i����@�|�Q�:Iz��ͭ�%W����@����J�]�
�g�B�fq����t��h����sK���%*Bz� (,��4q�sG��o�*�	[���[s@�ay�����HJ����Y�=�6}�NQ�1b��)KU5��[�1k� ۰���r�������9�k1�|էD��Bq��ɏ��֓Ѹou�w����D�VW�­	N��4ka��ϕ����YhH�F�q�"M'�8���m�AP��g��ÁB��nRRr�q�g�Ѱ_e£w�Z]�U%c��t�$ �Qo��w.�X������7�Βf�Z�L�:��u�vt�jT4��kUn��P�n��X�z"������?x�Ů���01u�����
2�aݫ�K��yP�ÅCz��� XÈB���u'Tĸ�1P����*P�0�6�]�q������f؝�7�f]t)QY3Pj�89,�"�o�0Q�L����/��9lJ*�1�(""o܆���N/�:�uGP�~�va����d�Ƹc�[�Y�����/�(_��]�M����Ċ��㯉���L�n�}��Ï���0�iU�X��sP9���k��U\{颗rV�(��o,0�<�������]���#�����Cֳ>mՂ]��3-m�3��NHg���4��9c�;��W�R	0��Oˮ��lUf�*��RUyɼ�E�N?��hPu�uƤޗW��O��X�S