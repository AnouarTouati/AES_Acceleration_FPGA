��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pם�Ǟ��(�WpS���<������	Q/���o]^�H��K� }��w���h-�c�:��S���p��Q%�W�q�&�E�TnU�ʹ�Nʕ�Ùn�y�q��h��D�`�<���S��,����j! ^��o�[}����A:��د.%eR8�a�6d7�Kg���p�M�:�����P�N��Uh�q�9M�nͦ�eg(,����x<:%G$����K��� B����ٿ�`TtK3��������̊���Ă!-�]Z�ę�*;��s)�D�c!��[�fAAj/<�%U���~b�v� W�/Px�y����u��m��_�=H��Nj7���B��@��ǖ�oFM�����&�X����q)��Jþy��q�,w����&�EЁ�x�ύ쌫_�Ʌ��2��N�4F�܏� �R��R�g�Tj� ��S��nN�K��r��������6�Hn��B�#.;<a��,='��n��.��= ����8=>z� ���2`e?�nw;@j��q�}�Z���;]�2I0Z�e��a�߻��K�Rk���i��4�(W��xiGTt.$��al�d{���� ����W�0O��P�$�0�#�
�^6� �r 갴�G�p��h4��V�ͷi��0�\m=����bj���z~�h/�9NRx���-ŉ�$DwB�
/�($��-�������#�ε�6!�\��<��:�� �|�P�T�� �[ᯙ�^��Vu�$$�967-$d8���OߊNtی������E܍y�s|_���:N/�?�M�RrP���xD-eX1�lO�xdhc/r��� �rl�O�bԉ��@%;eL�׉�e�*ګ���t׏ȕژ�"o�P屾��RB�?��pq�jYЯ�j�B��4�eUe5}�Є�J%�Wx��N?<�8&�C�`�o���ZB�G(8�}�d�yE��'��q���#����+�y5��KJ�i�ܛ�J��2���/B�M-��j�zvZ�PI"��$lY���7Y%��?�8�ʠ���/�6'#G�(Ż�U�N����|+Λ2$ۃN*�9J�JE������q=��/^KW)*z��Q(�
�R�8J�j�F��l�f����u�
S���ϖ��f`�0��k������\L���!�q0IE�R0:"b�1z������M-�cP���n~=�V�A-���S�����\�9���
�i>	s�e9s5��S��4<�$�Z)K�-���4����[E�y��vle����+�h�O�:5���R7T�
S2���ᑵ,'���^����x>R�0
{\�Y����8'�JGh��2�w?�����k$�g6��v��������t�Yui�������d��8;Μq�`%�O�^�	����%����瀆�-kEfwy/�i�d�Q�+�3��ؤ�8t����H������v"_��!�^n�<'�G��V|&z%�7(U ��v�3���D�$�l��s�X��;��*��8�E�Ǝb��X�j�8��I7t7_��/*]���w��8q�F���h��\�[Hy��^ܥ�!g(&e}����Qf�\�^l���?�O�5�]��5W���+u#a��xc�#⻇�/�;R�t�׉���c׃6u���YNh_��M�ޟ���h�ŏ����/`�v���?�W��ڦ�X�M6��(��Ql�f���b��1n����>�$�ƒ[jr�ތ�Ԙ�����8�3.����L �Ճ��ٚ�=YB�l�b���{s�;Ƚ��#��^JlW9����4,�R��`߸r�l,CO[l��46��"�{[��chfɋ���=��z�!��,j����.L4j�JУ_�q~������"��,�~�d��Q��ztZmO
��jG�Ф �c[RLx-�hc�GxY`� #�}��u$�����a����@��0�hY~��&�}UƄ$&{���A؍��'$�=��D%Z��@b����i�8��Ou_�Y��v<�~�Kc}?ܕ�U����zv�̻�9��]��Kp^X{.]��ߒS�pBx�ޯ��V��Nl�_;����]�����}�	�j��}©�ܡ�'�׷�C;eZ�x����t�s�p��U����/F�5)�D@�y8�a��$H����2iL��j�W�`�I�F7�x!�U�V_��y�(��䠠���!�����׀���Y�k����W/�Q��R䂅��;�x��HJEf�q�_�3(�f��p|�HԕB�m8Z5�LT���@�p�hR�����g�'��TH�cL'i�I#�hˣ�jc�#�(@��K�R�4�3�>���w�����ό"�	&9o2
`*=֥�xA�CzU�:�"��<��a���&3�G�w(���U��\��M�yz��"P���P�tq�4��Ⱥs�Q�������1t2��wKb�m��y�B^.�����k�<�Q�u&"�eQ�!�V2V�Kf��A>�7h$
9���X�4^�+*��N���]�v����`�n����6}��0��uTԑ���*����#t��=�T���^H��? �5��=4F�!�z��tt7jUMI����Ы�g���mθn(RUF,.]��׀��V�O+v��괱�,y�gF�2z�0�P�"'�պ�#^�g3tm��i���cD��h ��$�B�}���hl�c�=��T�:��x�AQ�=��rM���kNHUٺ�j��̄�&Me�B �e������HA��GbQc�4d�;���Q��Ԛ�8�;,�pTp��]�9���tl��.��2������<�����1�؉\_��H�q�M��,�ą���?X�zR�{�a"X��Z�C7����r���|�9�|w����iP߯h!,>�����ڤyӿOr<�E��&ݑ�'݈҅\���&�1r~�.�|!�.-�	�]�� ﯣ.�//�M?��=���4����4Q�����⏿�@��H�ג��U���������0��K��N��^s��S�[RE:��PKf�#��X�*2fȟss��A"S	=�q�ҍ .�Z�qc}I�C��~��zo`�S�"�)s*������O�`��x���#���S������O�Ώ��m����=�.e����H/1�)��t�(m������SZ�4�X㻍�O[2�f�es�L�1��(x���N�;Ko���Q(Q�WP�Ǉ���Y�6����~]��O���ڍTJ	˪��0�@�)x�Fu8^G��'��:�wo���԰buh/����l��2}��C@�<��A�zԈ��в����"E����+ЄJɇ�θ)z�X��6sA#�5�ZY,5��Y���o�c�9Naff�_;��G�<�Ɠ���d�mJ���X]�`5�4=���� �b$rY<f�����*�(+Ќ�u
�q��)���/eZ���Z?���k�i�"����$\:f���TT������w0?.�2=�Q�i���𺸟U��7�q�2�%������%�=��E�k4�\�ːg�OɁ�I�e4;۝�+%x����vC4��b����ͣNI��sCP'�VT,�QE��@�D$:�+\���p�=%.j�f�0��9+�/��q��*Uz-k����I8����>�4�bi�aSO{�0��	��g<��wgf��ZTc����P�x_��b;�ٹ�I�~괓rF��5UNjt�.�FW0�%�o�ԏ 2/�ɑ�����F�<y���z�3�B��e������E���Ys����ʭTd G��L�O��~N�ߪ�j�o$w�W'����c�Ԯc���{$_ �]���H}��`�AE棝ޖ�=[�M���	h�C_Ŧ���ۜX-�1�k$%��%3 y����q�?Wc�x2��[Ѹ��}����7���q�]&�S����>l�р�+=C�KH�M�mH �g�B��G8?�@�Wz�3�FzT����&��`�t;�<e���T�W�ů�d��z�𨫲QY��,%9B�;�nT�,���~����UU��]�":H���ybz�_��a���`��uȂ$)~��aѤu�%����9M��%!�g�p�RMMn�,��&0�Ԓ!Q��c�� v�ãL�R��������#�}"�,���rP��&(6���'V;�ͻ��[����Fu�"���e,4���B�Pz-C���$��W��ӊ��&��כ3 �<$�v�3���.ҩ�B�CT�A��LK�� \
�c߅�	pQf�1z��d��Pհ嬌�m,$����[`��3R�
��-Kt`8Asΰ��;�X�H�:a_��������b�x���2N�G��S�3f�]d5�+��>S����Pm:�vk樤�\��̈́5�/�5�N+'��3���[e�W��2�ɕ�y��[�?g� rK�#DpL���yaR.^�x�ָ�&���fX��Hf�Rh����{���	4�`7W�����^D���^�\���11%ѧ�F6{TGjk@���ma�6&@ܦY7�0��?V��k�?��9d����{�8Y�eR45��оP�<�
oO.`�#�W�,B\��ɠ�_�DkSo���)��,9����w�W��6x���{�|W�
�]��+��}ĕ�P&��-w�	h��!{�l�D���OZ������+�8��P .	I�Ɯ=ĭi��ՃS�h@��M��e3�!�s�#��,����b�f�Z˰�#��Ϋhi�v D�k�|�pfO.(t�U�֛|������Լz�5ZR�����&ց�!��(6�����M�#��'��$�O�ĵ�)��0.m7��*[��n��3���)J��}aω���h�K>��G=�%'���I�ִ�ẚ��Н|0+�U6�~8f��A���Th�$�W�D�eq���bB�;�PAڪ�<]\�-�B�����L�涩R���J�=c�P�<5�W
O�8¶S_��+U(��rYboA�ej�歒��E4$�OoD��N�ZT�Dٙ�Zys��9X\�����c�"������. ���GE��p����ߜezgbFiө�*��l�c�PMX��ӂ;L�B}X����~�C��z��i]Q�np[~T{}�-^=ݰ�@���qs�m��{�uq�%��@vM�&?"�P��l�wD��ӮLWi��FA�(�e�P�HQq�����3��Ӭr$;���'s�ߚ�T��}� ��O��[�O�-:6��\L6e	ϋU��TO��(_]�����N��,�K�<��L&��8�4'h|n<���ú�@��:�RL���z�ɽˊ�kc
/��Gq�Ot�8�OH�s��._�	����~�]��<���rTGGS]|��uR��	�B�@a��;DE;K���޹�����*_�hҽ�{2��}P|�ƇO�:BH)���(˧�FbWǝ�q���΍}�T%m�G.X����0���a@�<�KG<;>�|���.�2��,�![������
�-
�γ�������y���H���#��V�.D�M�?�&��q��ƣ|M>���­�-(E��_
�~P�^�X��*����񃶨�y,1�B�s	���X*k@x�&��c�kWF�/�����us�a�A�h��,,n����<S�����C������u: F>�@(0���,�����p�*�Ͷ:����T�Fu�ګ�p�=|a<i�a�p�MmS]+�FxG_��}2��;B�u���]��G�uژ���?b���h�k�"�f����?��xRb
�W��ٞ_*��<��oZ��/�g�?'�QO]�n
�B�y	�? �N'>�pթ����1�,�N�]��tICk]�?���Ҏ�_��f����p���9#W:w���	��e��"�=���'0MȦQ�_?���P�g",K�UL�Yv���?'���#Ϳ�K�	cñ=���Z���q`�>PT��nO��A�dqM�g��Q��� 4sѫ�w����<&��k����	���7u;?U�x���w��`���5� A�x���a�+�H�採��b�,PG��/��B��f�7j��Ğz��[`ȳ����').����A���w#��i(/Z��~�DL��8݉
t{ 9�)�̢`��|��W�pT͗����bfUhm��B�����EX�fis{�B��Hp�����Ӝ^bѤK�i ��W1W,O�M�C7E8tTI���3q�}�TN������q(`�]x���ѩRNQ(�kݾ�u[&45��vB��Q�%d��Ћt������n�(� C1��Y<�?+&�,��F�IG���%��IՖ�ѡ�Ӟ�wH]�ϊSl>�<R��=ݨ�W�T����j\�%e+@�%
4%Ӌ����'�f%כ��
�J��7�LĴ�"����<�(ǣ����^�_|^�@��M��mP?o�%�N���h���EۙA�)f�:����Y���� �V��� �Oy����P )ߏ̡��l��"35ڱ�
U']!�)U;���E��Y�< t��E��.�|����޻����`� yQӽ�^J^���n|�!-ׅ�>���ЇV��܁�8{�N(�{	��R�?�Q��~4���e�1��t"��<�_¥E-{�B}G��r���drg��Xa;S���$�V��-z��W��:�B��L�0���JR<S��o�I},~]uαD��q7�t;9�B0�\ܹl
u��!G�5t�Q�TM	(S�z��:��ب�'��_�=R_rJE/�$�����t��iD�s��G��@�0ju��k
2�d
9��{������YW����+�&S�ޞ��/�%(�A:P�EW�e`-�-is�N��	�d.F��=���me�K?����_�I�\��%�"�*�1��Oy7}�p��G��� ��w��w�7�-]7�j����g�=����Fxտ�	s�}IZ��`�<ϥ>�&�� �Kt?	pΉ��'��~���$yP�x+a�����n��I�!Sa8p����P���j@D�Dr������G~v�,��O���3�v���Qx2$X�ʫȔ��q�4��ؠG>]���U�����e��iW�e��+��R1%�L�F��m��2*o����������_������� ؑ�{xú9]U�Q�{����HP*DJ&$"l��#��|v���]�[3~*a{��h�uG@0�@rIB�����CR)��E������]��BT��m�_R�K����5��"�~��KT!�� ��I��;a�@<�X�V�u���v�C�[���sX}����w��ҟa���B� ���n�+(3q
����UtG+�L��7�hs���S��4YZ�Ԃl�5�J��;��P�Rv�j���'�U�U��F����d�K������}K��X������h���n�:c���#FIu���tԋU=~[۩1'�U  2m$���[��'��i�s��W=i]!�a����u�����F� �&�P�ݸ��h6)��I{^D�r7Y�{1J�V[�͂��ii��0"{�V����ۡ�}��I0<�O
7}��Y��u�C�(�C��#�P��d!%�V��Jo�]�����P�bm�[)IS�W���P&��ȟ�i��m��Bb~B��m�r�P�閤4�B�ŕ'�G��c}�^�<v*�f��T�1�_�F萤y9�D=�:	=���)�0�-���ԎHb�����r��zr��)Vh��_��֬e�5�%�����+1�B6,
9���y�*d�=Q�"%2���I;���|��X��Wkف���hh�l�ui�*��=�M"������Q��J\�%Q��������� �%�X���u���W��߼S^)�u�^V�$=n�P�O�"�`�(���E'a�f I���t\�>��%�����̖��ʗ�s���-Y��/�S��5t�MA�\zb���=�����j<x���K�w���@�e~M	�h�pe4�~i�RyI��?	�v%��TJ�tͧ*�;nd�0{3����X��p3�VhDa�xX*���Pu�T
$�����8�Y��ýo������T7�X!9�ەDw�)������ Q�U9������R����,�Ji_Q�l�sY|�|����9����P,=D�]"��T�&	z�8�K�;�����}��a15��®�����H���[UAW��i�:c 9�o�)� �e���� K#�w��v��K�w�����&L�	*Zz\g%#6ѧT(Q���vl/�o�/�4>�.lY�Iyhg��o�0j�@ϗWbN<x�8G��lh c,LQ���G��uW�R�.������_�*������=�-l���D�Fg��\ųh*9t��eO�b�uͽ�f�ї�&�[�'w�{bŐ�>+Yt\����r�df���5��".G"�Yu_X<繈*Y�e�iZo��c�Ssl�
vӋ�v�h����j�G�`u�Ť�+ XF�Z.���s���|s7��44Te�[�������T*�&�8p��k����cD�'!��ȉF��SǢݧ�S��	F�����@��('�?FtG��:���ޑK����<�\K§&�J�&���j��7ztM���n�v��xy|�xT��?�w������b�.a_���=�Z�E��LjV�e��I���8#H��(�o��������`�H홵�Ͻ����!�=fa*"Ʈ�7����qt(v[�՟��J���N<T9�U"#+os�{�����),����⑘�ʉ;75�~6���B����V8�X{��,�ȸ>�g����
����Q⭵����ň�&~
4�؞����cj�-�ԇ����3'	8����S�Cy!�OVݧ�W��Nf�!%���x��a\�v��W9�y��0�c�/7*'!]5)7
�%}z���E�|B*H^��Y����Mtᡞ\.8��N�^0{�@k~H�ʢdR��ю��1�(e{���V����g�ˁ�/{k7�2	 9���8�ѷ������uB\S�?$ F1pN�~4k͊C������z�'U� ' p�_���9�@xq�ߺ��~glF�������u��Ìx�uYZ�>��5�iW6�Ȅ�2<l��X��)�0^9O�k��S�L���h|�P��SSU��U�X9�����u#�
���-�bNB�j�BfR4N�b�P)�,CM-�՗��՘�`�|1�j��"���;3�<[�E5��2�-���B\Sa2�q��	�ѥ�o���k�p�BB3JڡJkh��1���b���8G�`o(��ߊ��	��֋ք)��#H�m��E�D�?8���<���<vѬ)~��U��i$K��_J�	k�)l��%�aoQ���ƒ"t���ǴvN���|���-�����0�֫Y�sL�E}�'�tt�r�Z�X�YgԹ���F@e���|Z[�d/&:�3cf<�usκLB"���7�0�~�A��J8{p	rx�QY�j��L7J�����įAJ ���hgQE�/<䂲�d�F�� ~<��i޺ᕲ*��>�C�LE�c�ބ�8�oazӫ��1�M��JpoùFJ�Hhk���⊞�M$UP���$��6l�/ă�$�4�8mv��h V���e>-����T�7���l��)����1c�2 �?U(���ѪkcD{�^�4`+�0W}��H"�;:S�3�B�Fȗ5^�!�׭k����U2
g"�t�K����6(	dc �o���
~����d;�o�]��b-���P��_�g��!�5l�v����:-�dg�2��}�0g��+N�^�Tos"%�ʹԳ����$� ��eɎ��Kf*�y����ʋ��Ə�?��ی'��6/)n;� �+��_���h�"h"A:y�ER��	;�{8Lon�3��U!��ń�Z�x�.k���S��ԋ��Cc�|�+?�v� �nvu�r)�k��v�h+�# M;u���ı�����4`������lz����̊�*�}��q�K�����,���?x픷ʿ% l�$`2D��,Ҁ�5�d-�)+����:���y1zI�7?�WJ?�l�-�a���¼=�h��#���9��d��^5��?i���o��I��������x�5|�$ЙZ-Yv˓)A�P�w�6�J"
Z>+�(�d���ö yS�X"ber�2+p�0�9h	��\Wab�	sk ���u� g-�&�$�:����;�6�x�#��.u��P��"yo�8ݭU���&�C��x�A��N�����t�J��۱�_Q��j�x�6|�������8Q�ӵ���|C�{�ңX��� U��m6�Lk���ͣ4�+h������wf�����{����C�b)r��iN1v�Jp�f��6W�F)���>��>�%�G��K"k� Lݿ?r���������Cx����F����J�Y���>x�BX�Tb�M'���0s�|kM\:�9��IĽ��讯�y�YnE�GZY*�fRK�:z���8�A�o��D1,��N�[��ŘA~�?Z����JY$���y���