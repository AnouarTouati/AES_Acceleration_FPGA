��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P��/�͢a�-� �9��@W-��ϴ��qd���O ���Q�#�PP�[x���
1��m΋�E����1H2ӑ�~�l�2�����ա஠��|@\��ʎ����/+.x�E�)�J��	��j�����
��=ϥ�X;����������N��]c](�w�o1���|��t3��o��%�`����`��f��qv)5���Y��S�`�$*�<?z!Z�x�X�ܾХJ�i$\)�'}ArŸ:o���C\y��튩SHo�W.r��(@r}�A�;�/�~��a$�D�}�4j���ؒD�߱ڤ�y�Ż�D<C�:=���PA_�|�2ڛGcD^X�\ߨ��_�SΣ,`�O)���Hp��[т��$���J[���WK�� ̀⺔� ����̏�#�`�k���)`�,��[�}�XybI�M����횆�ga$�vyЭ��[E�2��~T�;�w�ᶙ27b�Y	+P�
w��!~\�Y2�����Xtp�P<f��n�����!$��3D���q4�,�0�4���zN�z<:�(���{t�e<�O4<�J�\kP&��h�#���z,�-��"��ԉ�z��.�)�&���mϙAJ3
ANL�;�I��q���R��[�rh��n Q��Ê�"ۯe\�UK����]�F��Q�Ea�M�vU����0�T��[��5h2ғ�ϝ�ώE6AD]�U���V&~�3C ��|��aQ���#�d��D5��ʒ-/��AM�9�8kl��ȥ��xs������\C� ��l'x}���h���E�)
>�gB�f��߳	��>(C����g[�xҪ�
�¯��60/���b���MÙn�+��F�:�����YO��>fY��sn�=x�R��ocj�L���G��Bi�[�z4�� V�ݫX��P�wj4�q���Yjm���1�uk�Uk	�`"�g4����~��������v�`JIXU�]P`W;g�[,���9�%�h���T�����#c���ßڦ�B�b�8#���`4����d����}�#��5M����*���szA�ĔXB��,��{`�z#iWw�t�k�V��=��-�0��ݐ%Lx�z��g6�l�x5���,+�+�ha�����͊Y������9�0�
GbhmAZ��TY�х�t�q�(@B�2'5� ���L��y@�2=�uPf�eHk96�����д����*�Ws��)|���`3o'�KAA�7;�YL����ɃQ�*�Z���i�ͩT����0�U�1΂�H.s��H֦�v�}��$+�Ď�����x:�ґ��ѐ$7+4WN�a�4F*ֳ�e���g��3f�_��� ��5>Y��PѷT0��Mf7�֋���蒪ײ�X�o-��֞b״�t�o��8�K��B�1��j�y�"��lzx̾���x)�P�^�N܁�bV�-�S����`5��$��TvA(6�����PA�c.4*ĳ�?��䗔�a��-%"8���}�tiu��u&.�6B�m�$�V���Q�8����MJ�[h1�f�a+����Qf����Е���ʎm��~`)�m��'B���E^��4�;k��x�k�up0�$��!��Vp����Յ���i�r`�,����C�(mG��f0�Od�4փ`�9\��\�|�r�wU�t�����H�����s�.�:�`9���/lb����CW�4�n�SQh��N�I'R���,_�hKu���!@Ϣ䄃d��n�GH*�ȳ��h��[�H���i�7!li��W ��5�Ou �	0��([ǆ�$p�F����~�1�<G��x�����a�?�����z=�r[���L�s۰0?"ٙ��):k�Q���^��ה8Ι��p�ܑ�e��-��M@���e.���L����
���(�\KG��P��<��f?o�8��`�ܔ��w��-J��2�`��8b�6|���<ʰ�� <���{����>L�E�d�E%�c�մTX�:�a���F��w��71���G�a�NX�5.=�<ڮA��~Rg��l+�l��.C��ɮH�l�	��V�Y7i�l?�� �z�5+`�t#���#�#��*��@�ʤ����2nD�����V�j?�:]IF�C�Q�L�ׅ��_N)gH�ԙ)�H4ʖBbEe��m'D?ELv:C�_c�cL�|ĸ�J�N c��k�1�l�#Qm'&b^i�4甐 ׀E&r���u�N�mf���*`D6�PZ�������lT+=e���[��� ,��x�#�O�,��Č�I
��ͼ��b�͸��h[�S׉0^��j!��r���t�l�4Ίԍ�s��0�{-���XD��{��q��)��BC�c$P^�kZ+x���e`o��%S'pq�l��;�f�S2z�+� �r����F��+v�D�g( ss��JTV?�e*��MY���)J�+�-p��I�Y���A���z'"D?X�"�$#�v4��	d��{���j��[MԥG�gJY��1�n�]O�u�	i@9���������y��(duN��_K
.
�M�����8|��5ό$4��:{���G��C�eH� ���e�=2�]4q!@����!��<�@m��G-G��Y}��=�������E���ˎ=`kn�zG��s��3�8WnY��s|F}Y$--��#x�tUkF<��&��0������O0��JDq����'_}���[k�!�c#?I���q����?'�4��&-@�@�1�4ٳ�'f��~�0.p���l@�:,�n��G�T�1����OH��"�������8i�R��Sà�$o���ze�F�C(�
��5�$
��_����@TS�����r�Fn_�UϿ\��ƅC�5L#Y%�`L OL�����/����<�C7|�E;���=fX�}��@����ݸ��2E��e��
іoį|���C�����_��,����6lC�d1^�Gc�@�����r!��!
n�$$����<�XL ��ku,�����EC9���z˨҄*<�I��{�뇇rcc�sXzK��]��`��*1OdUj:�W{��F>MJ�+;@O+;��B*�Qt��[ Uz��f��4%%q�m�b��B��j�am���!��;1���5�(��zX�L�� =؎�Q|�~eȜ������e9��4&÷�>��l��`��L�ټ��C�e����V�g�K^��)�� d����,��.c'���KtheD"2�b��9l=����B�^�A�ܢ0��K����Q����߾��{_��PNU���<�7�s���UX�����L������S>I�ą̅`�� �Hӣb"���������	�����	c����4�)��x��kO}[�� h<ө���'�;k���Y�Y��kZ��rJ�}L��Z}#�~��K:%`KF����&���j7�B�����F<z
��N������q&�ߋ*�>��f������|�4=G��D˘IJU���R��n�9�E�������H/��TRn�J8�It�\���[�]�n"L�k��4�B��
@���\5����tG�C.� ]�@�~���I�yv���]Jbҵ�h_ـy�q��%��aA�Y�tIـ�Q�g$�L?�,�����ܸh4���X71KF�Ck4�׀�T�׼�/�.^Iw��G�#x6�?���?��#�H���if��U�Z�{����#�%��E5���ܜ5�9���� ��y'8�J��WqP��o�魂��m2G�B��x�N+�*��BJ��4��9:W�b��%-=P�	j�La�|���,�W���{�^��
����]ձ��`��L��y����3k��i�p 8����IK�8\�*��o�Zr��}����q���4�� 0���N��b.LM�������Y��Ȭp2+K%��%�{�4]Р�X�Ż�q=/=�'G�Ϫ�a:ݟ��y�o���财3�x(&�.!�,5��ʷ��n��������fB4!p�#����\�KԬKh��DN�Ǌgp�B*$�2�D�� �(��.�+@ e �jd۞c��T�.�sM��F�8�����P���|��@˶��xS����ޣ�2�g  ETf��� Қ���+1k5��>�Ų!��g�w���kEn���ܥ�J�/�+�k;J�]3Ls�����\u�W7Q�c..�ky����U!]d�ğ�C�g����������'���d\g���&b>h�	���BX�!�8�/�Y��@�\�VymƁb����@�Vx+�Mm]Y�oX�oCB�A�h,*沈>��.Q���w
wvh���_��Y��,��~��x��]XBYz��Wmm�}.ɚ�k�~��j8�����Hj�睿hY��7�ݭ21	��İ����e���~����kY�t��g(�Ţ�?g}���>���ڿ����T��F��\ݎ��֟�%!������=]��Z��t��P�2����'j��ӚW ���N��#Nt�4X2N��O(L�B��^&%�6�m,�J�v�f��n����VJ͡����������ri]��.�}K�X�~�	m��k�߮^�qa�{SΚ��ʺ�uLV�68j�j� ���T%Y�L�	f��q�h^*Q���r�T��=�XaW��<ן���ljl����i?C�Y�>��E�^�dk�w֜k��Uw������#]YJ�ߗ����MА��3.L���i�@��Q�p����`Ǖ �����D�1"M�ԝ�~Ȣ�*����<TQ�5���O��~oO�,��jtO���~�K����L�9�����l�&����J��t��7ԒP�3���s�x�%̜�m���͵Ҷ���a�i��	�f�b,������;/��1�o �t�ޘ�c�з�<�=wt�y�A�Vf9�I��BW�A�]�}�����)
W��1f<�*�'�PE!?��ϴ=�j�G�|�܈���K-�z�AD��a��O�/i��g#_��T��
[�j���Ʋt.��oQᮁ�t���ɛ��1��(Jv)��+k�G�剛� [:&ЧS{+�� �\��<$�/��a����J%��@?ſܷ`��&Ɍb�q�C��P��%��zp��r]���KΓ����(iv�bp�M~��$�?�9e�5�7M�^��ml����?�1��Nx��,�n9�'V-��4q�ؔ�M�?S�ɿ�&�c���c��S����)�N'a��̔J�G>��%{@&l��A�a�;��H原x�`�RP'����rZwh�!�Vhb�qS V
�����."��(|��O4Aaꠀ Za����;K�X�H���w�g|��
�Î�x�.zwL�W'NZ�	��v3���R!������lB�c���N1�_߶LeHmS�C>�Ƙ��Ɛ{�Q�aRz5`���%���7?�b�Q1�N�">��O�g,H�_�������+��-�'�`O|�ݎՇ��쓘Yd�$�2��W8ń)�
s��H3�?G[w�+�\��	{�	s,�y�g5ʱTS��(�Jr4����fit( ������'�@�w>:2�"�.��1�V�Td��ͽ2�ʻ$���V$�r��$�t94҄S��!�8��}F#ނ+le9����C�
p|W-��
�f�.��"O$�5����"��� Zůkn�fP)hA��>��9������g��DG7AB��A��s�����%��,�b|��B��<�2��@m���τ5��u�3�Ҡu����.u9�*=������R(k�ƻ^5	��3�?������جES�W��?����@�@�v��RE�R�0�-��ļt�����(p���[��estS)��,����T8E[���MT�XQ±�F���ٰ�Z ��t����]D�$���a�|���U��LQ_M��y��q�[`�Y'��v�v�{�"��X0��Mq�m�E=�rY[����:^w��ЊybY�h�`�h��&�@��]=�ޣ�Zp{R<��7nI��F��n۬�G]��)�@�%�TL<4�>��ܖR��`4�g���ԓ���4Yě~��x���*~K!�݉Ls�k9כ-#�w1������u�2�.~��q�c���6Uv��V���h����|��X1�l������/ �K���b�W�)^tr���ʡ��'�r~�WL[�Z��&Q��e�H��9J��ɳ���.^�--���'mSvA>�tt��؁��b	c��E���6��O�sA��Lw�b�0����y�����!״) ~�? lPD[��15(��V7f�~�$璭���gw�3�7�Fw�80o���n�/٪U��K�)c�qJ����2��h�׊A"Ț���[M�@F��C�:��Wx�y����;������$��gj��a$����%�I�1ݸ���Oi�˷������n�.z�W9�X�Z%��[B�7�,��k�h��1�ED�t �R� ��Vj�3(��֩�
������]H�Ic�$�g�dW���Fk}�2��I�J�5wTg�(�:D��?�S{�����8
���s.Vr6�wl���	P[��0w�hĞ�K��R���"gr�ҙ�i�����u���@��Nl'Ny��х��ä���;���՘��aW[�5�0�@M'P������:�*t`5������V�`�Ջ����XR�$������W�jrj9κ=��񻒋�5���̿�K,���3X[}���֬�����Rw��!C�m�a�ӆ`�i��(�Tk)D�t7ӛ�#irP�y��$��``E�� ��W�Mq�\DZpp�%�7�G�lE��ͥ�X�7�=.�MU7m+�ҁǓ3A�`W����V�����II�;(���!��v[ͫ��n�W����D��?�)�e���`����S1�~P����r#Ɗ�S��7ⷱ�X\%�M9�)[f�]���؟_V�145��U�0~�`1�T���5.r�Tŭx�1�@�Gptxr��K�5�{V!57+Xr�H��a���[�9�3�+�����x�J�L�hQy45�������-?0j���h��ܟ���8�4���&' zJ��y_�������=W�ѹ��÷�)G��8���`'�"h�gUr�UG�a�h	j���@|���vL;D?*������7���|��lđ:{B�޽��R���&M������\~�* ���K_�hi�nk���><%��s��wK\��h�2���@"1,�@� m��ŀ.���.]��Lb����lO��zDD��O�w���M�x>���Ùd�me���A2U�߰�K���M�} ~��.���.����l�X��:��Yb����G�Mvq�����\7J�l@Q�͠��+Z�!�/��R���т�(�� �a�
����ۢ�E����~����+��0~��?��
X��؎�傶
�<��{e_�Ҷ�Zʤ��۱�[���>���>s-折�sX�^�b��SnRj��1�=L�{�\ҍ�a���"Y�@�tcd�������Y�0�?��Ћ�ť�h��; �f��=[uΩa�f����#�R��Yx��s����~��z�\v��Ў�n�H듗��IS��}߂�n��[�Q�us\��PI�W����<B�
�Q�"41'��<��И����G��u�.�9�����@a�޴ɮ��ɣ��γC�g�R�A�R;���	�/�@B�i���/�a�f���Ys!�{^��f����{̵�@m��CYNg��b��utٹa�P���шj�ld�=E�4'W�.�Q9K�����o���c5�!�"q��TL�I�����/g���H�`�����1e��Jc�F=�yY+���L�ɠ��m0Bg�'��?Ap�3t/�B�,�r85�`7�a{���c�Y��������B��wnO~�E����^�k������/1BM��z9���[o^���U8�� jK�Bj,K�1�P$K��L��P��ўE>>s��&�7$+���~̓5�Q�6&i�2�I4�\�D,Z�o�a�K\p�5�:�qдH�N�$Y����r��0쒌��\x�Ay����3Ԭ����;��6d�n�K�I1o�J��#�6m���۪a�o�6\������Tߋ�F)Z,T�[PXW�I���D�6s �~�DH�uͲ�lB��$a����R)�1�R��{ÄF;dD`SrK�j�[-=*��1;�絥 &)R#��H��ཉ��\�)��-���O�l�s2h&P+����-�����$����;��r3����6_���VK��]Gm������H�7K��6�:�B���Ѹo2hM�4��6U���}E�lx����N�z�(g�R[�C;z�ia�;�������"��THz}x��0^%935��;�<W.�*��󰪧M�^[���K7X�3IZ�j�ل[{W�.�H����E�i��o�:"y�Gl^ �SF�A��%nD��-DW�>�b��5�u����;WKs(�elf�%K�0WaI0
n���(���3[e)˩o���Ԧ��L�@��C��'���Zܢ��
�@	7<c�ok]����jȴ=�U�H��E)Ԍ�X�amj���4�"��Ċ���v�h�Z��@���x��,��4T�3���q�&,��h��OFe���`:�.��X?�K����<���؊58}tm��@��M'D���V���9�P3ݮ[Mp�틝?�]֫�.�/B�'����k���`�SL��v�Ż8~�����+r��@$q*��O�v�ڔXB����~�a�W��F�t.��#��yk��(�<i��30�۔��R�pM��k��C��t��.L�1����E}�+<��p�������d��$��nz3U�����v:���p��W%@�u,�6?j�L������K'�޼�'X�����ֺ��iVo뗑��b�ʟ��7q}��7Γ�8��!����2�z%���3>2���+�8�{�(��`�ȣ�w���N�s���9 K����}�C<���	�$�S���g�1��}@O �V�*x%��^�Sp;5�Ց�5���P,B5w:�Y,{}�N�$pW��Es_��p�R#��޷�$U��-6�d�רݨ,UZ����W8�zl�4�L��\�ٻO`<��{�75>ģ�����L��@�����׌��+Ӏx��X�+�//�Ŋ�ٴ�x��ƭ.��-#��%}=�%84S`�Zr�������0�)�m�p Gh��TpQX����[�j�s?��v��%H�B|��� }g�+��
�>���H�i�]3��������o`%`�D2��i�c�a�RX�Hds���}��
��)	C`Z�F*
�_~�c����Sf_��	Sm�����>��db�k��$���B�^����\+(�;¤�R�#Ss��S@���ݱ�P����5��-�i�u)��%W&��O��Q��nz�b�"L�i�%ȼ�L��̧%��yHc�},+P���M�^J*��s*D�����&R�޵p5fA�+�?�%��d�F��o��<�W�q,��n�탫'p(x��=-嫍��Y62a����c f;�Kֆ�����1��{cG�3aR�'�R�چ�瑏`uXt*+Q��BX;n� ۅ�Ë�I��~71;x�ؼB��Z�z:��[�w�0!�Ի��Pv�.�U{ؘT_MJğ�kEPA�D+|W��BU�҉���� �h���Y抙}WIa��?9�h�kJ��v��ğF۩a��!35:�dU��w�&�'�D�{�փ'd 3;_�[����4�b�A�k��q���5��LѠ��5�Q�&�`S�B/o�#l3VL�Y�v�ZRT�jr�3O�Xg2�)V:�<M�K��҆ �)Y?�`��ܓ�Q,����,��^�X(��Յi6w�'���K���H�U�Õ-GߚU��Fu��L�3���۪ɛ���r ���*��k���M�>����k%�ˌS,�`�BL�&��Pc���;U������`��B�	��ԍչ��$cI���)��crL��ub�(SN}�6��KH��x�G����)̈́g�]�sk��0�'2r-�S�d:K<�@�J��j}��D�\;8�B@	��������e�q`6�K�?�=�jss *4T�GR����ci�D����2�U�P����U�Ew��N�B!��V!$[�QS+�Χ��וt�] FR�V.�k���	.+��5��WC��5��>�6��݅��|��E��f X2�]�)ҶP&��v�I���j�<�xȽi���>��;�5@�G��LS�F�]��H���/�m�6�ޭm�p��ɱ6�RaI3Uo��veA�v���$i�n��[�zH,���k�eM�P����%�şa��|PC8� �-��~��t��e������>	ce��.`����򸽂��s���Q��&��ԥ�o�]�'(�B���QeZv,,}/�q��;�c'�Ŧ���sKo?	����x��!��4���Ln
k��:r�ດ�1/�����%�r" �ԧ������Ww_R�7}���f"|LRgB�f�!�ӶÓDK
_�
�K
�Fte��e�Xڿ7�@T+N�t*�����ފA[�v�`�=�ӫm���h����;�7�a�A9�l����82�4���)Ph����9>���G���V��ic����G�Z_����t�׸o&Ɍs�����Uf&R4n�^;��8BW+�����A(Y?8ɕ}+l�af[&:���~m�gW�xotl����<^B#�xsV��\�����&�㙒�/�N�m�Tļ"�Kc6�:�dc3��L�X⭙���U���v����p:��A�����w��p�"��w1���V�j������F��U���s�v�:����5�o�X�K�B�:�I ��pS�q�2��?R��O�#�Ϩ�1M�ƀL0YD� ��l��N�v����tY�.�C �=�
dRy:�����]�:>��p��"�O�B�^X�fd��b��^��˒\2�m(�����Va��ր^=�m��/��&u����bA�����@t�9A�2�Hd�]��+ H�*�}��m�<{�:ٹ~v��'P�l�*�3���]�:Y�I�bk�����[[��:�د��j����>�����RR�cSR��atż�?������$!ac�(���������|���Ֆ �����-��G�e���.	Y��0��g3�U��sQg�t�O�^��1�4q5A>^��S͜�O�f@��D�Gwj�b�˺?c�=�ӥ�q��K�В{��jn����7�n?9qkE�v�l��K���/i(^�af�X�+'N�F��(�
��m1R��BBv�p5PI:�$��K$�Յ���7cp�7z�]��w�+�����i�z�,���s����IↃ��ei�~$��XmN�=��il\�P F�ZR�n";����]DW�����K�5pjȈ�������� �$�u.��G���']���ڱ}d�=+���r��}G�9�����b�tUl�V|��?��,�M���x7�o	��Y���3@?�ā,~�3bN�l��nc73���8�d2��Yn��d�����3a�p.:�z~�rA��Ŭ@�ckpx� 23O����`I�ԗjU<-|���_�q�M4��	��L��Ց��ʵ�"����dy#k6?`�u��X��8q2R��~?p\{}TK�c���!U]�;7�	��5���Q�\�O4�ٔ�дa�?B��p&O%S]��P�gL�D�I �v��0�,+�GV.ʡ@� ��eO^)�v�H�n#����
�3�&}��r ���x�,�(���i!�O�����9��j�P�
E�
M5��݋: ���z6�����O�֢��t���]��ܺh:ݴ��/������X>ټG^�c�Wd-����
���h*`�L�+�ek�x���g��!0��)�qH�N�+G����8�������f�����@7���,��"O����B1#�Bl�%��D�F�A�Ymv,�.�ՓA+���%�rOc>8�B��`%�ȳiF�*G�� ��k��f5�Pc�5���pI�:4�����}��,�j�������Cp�s�MI;�����D
���=�ӛ�#�j�>�<MC�+y�pd��2��o�p��-�38�."�[���F���ZF��e�t�:/6��z�f�9�յ߾��|�H�f������T�p� ��B�Q��V�6�5��<��(-}��c)r��aW�~���kk�Tnl�r�ܳ����8�����j,vg�R�x�c]��*r-ӷQf�Pʼ�IfM��@�%N5�Ŵ��?Id��Q�N�G9�x�UG���n��$�n�/�
���Y����#�r�%�h~��l���#g�V}T�y39s:es�����Φ��;�R8Q�	���v��Ā½�"�������|E��Y�~���q��\���=��.!�0S����&���/�^��LD����M�VL[ya�m5�s:;����Ѿ�YS�\�K�/e;/;�-(�t��ͻ��ƚ�K�Ek-)e�9+�i@����[p!8U�a�`&$��Uz��ʑ�+��s[���j|ۗ?�!�S�=�יsw��u~!��w�br* �mŠƊҚ�eE �, ���frz-��A&L�P��9_/Ю��oS.Ǯ�=U�؅c���U��\���]`s���o�MY�֨r@jWY�>.|k~��zj��խ�bN` \/����O
LJH7�E�c����$F	}����|"���~r
�?��BkAy��f5�E��SS��7QD>�G���3�j$T	�Җ��#ؼ��t�A�[E����_���0tk6�Z���M�ӑ��aB�	+������X"�q �O<��FIp���nR�Zy?�~���	�ʆ�OLΟCn}c )�L��I?0�U��Zv(���#1#�8��5`dԌ��a�v��'�8��lܿf�SP%�M?
X�����	6Ҽ����?��b��YY6����g�I�Rny��2�<��ڼ������	����OFR/�����f��P���G�Ja�kZ�a�q!_>ᇃE�r-����Y[ԁr:����}Y�2�vk������(�J�y3��tP(������2�ʄ����K��/+��q�ZMO��~�\��9w�����R�wA�� 9?���x���j�A{_7K}NT���d�k�� ;�W�azS�e:;������x�& ���T�aX���|�1��l�^�
'~%�[S�T,6���t�΄ɭT.&���~O�F�x+o(0i�
��@D���,���jTϷ�ۗ�Yn�����e� +O���?cݸ�b��ƓR�ѝֲ������䐣o��Ң��M�a��F'�󻋺@���Xa�z2[�w׍�롖�㏰
'&M��V�/�����f	��/�L"(-�E n�*��Z�������fr����]8vIj�N��X�
�59�\5-������mŠCZ��C��=B����a�"���}|���#����N�w !��3
pg�[�����B����h�܅zچf��s=Tm�x�2�|�q��K6�K�������� Z��[`�^f0D}G.�	O2�F�*9~��"�6�zuS\MT�h���_�BRA��?���`i^���=?h�⁯����W��f���`��"�t #;��`m��I��"�#��WN�I�L,��-B�-<C�-Cgj��+���p�q$&�^*�Ԍ��#ǘ��n,n�R�]2Κ��.&zͨ��-N7{��k���`���ݰ��:;���S�-�q]��^�Ix_��hU��S+���ī K���,�N��ϻ��c�(�\mџK#;�.��X�� ���38W�##QkN�l���];���6������c��[��v��xUՀȴj�;`�R�\��Q�|,��u�fK*%t_v<y�Ά���v1-��G���j��u
��,��W�Գ$�?�!|�6�6�D<n�}�����j�P����qu'G�C��ι�%I�g}���Ir��4T}��TKԐ.��{d�ִ�w%:����A.g�����V�BG�YP�Ɣ���L��aѧ�3W6�t^*�SQ��xS���������P��`SYV��_��L�?��ڥhc�%�I�][ok��H��X0�L�N_��]�6�{C�]P���!Y%r�W}����]ET�:H�!�K�YpN燍d���6 !aS<��Q�yAԵ����]X'�rҘ�a&#8�iT����Z?��N6ꥠ9r1sor�o7��x�3�+L�6���L%�a��d�������"�Z�>���XN	7��Zj��=9��A"�쒑�
�ªkӲ]���>�z���p�\[NfGl{m��y��`!ʦ�s�jk�{mew�RR?�z���T�M�/o�����>B��&��t����;��R�A!��2H�)���*�E�Ɣ�>�6	�Q	j#҇�m���J,#�ʦ)���r((�M:���I�=�J�y�;k��c���n��匼�7g��:�!�-�T�:6i�[	��\�Jb\X<����[v���!�c.�]��|����̛o��Õ�`��5��{]O�w���b)���=�Ք���XA`	R8^�2$d�Ѡrr�9m�uC{ט_a���t������$随�_g0�വIJ_�X����S�>.RS$���dy��-����D�,�]8*���M�s޼�g�<s�2��l9#�gpH�x��ߚ��M'�K�8lXng-쌤XF�[覯p�ho�Y���$���ԿU�n��F�����N�8@��5��7|d-Uc��T�'�\��.��� rKO�}�CR!%�l�1á^���R�0_#�����bTX�� �n5��t�NJe���D�j��7���;��뎺J[4{`�/� 9T8��N����r[16��d�N%})�N��?�kq͸�w�#))?��9��iŸ��m�*�xǳ/N7<h@T��J�}�j?J��(QAY��Z���Q���r�n�jL�8{{�˞��^����\��zio�R�0ئ6L�B	yg{Kg�Ci� ��~oFL�$J�������9����KW"�Bv_��z@�F�^F3I?5'TSG���|��Iի���8���%��V���1��VR�>$Ә��f���v5��OLrbz$j��Ey�C�8�K�D�_8gA�Z��^�����0�i����=���_�������Yq�m����4�4>NL�.*�j8i��@%�DA{�Cjd�|��
����̇ք�V%L���f�"s��R������b���6�	_�pq����ٗ)f���!]n���k v`(��'O�8��È�O
R	���ﱯ�xzH�k}��W�pL�����&pP���J�<��z�H���&�<�L�"�ȍ[�"������C��5>�:_�0',.��-�1�z���7o%�/��������TD�J�r��?�F��6	׮���!��<tew������H[����c�` &޿c ��WAD`:7W_��Z���4���["x| �4;q�t���5�;~�|�v��NQ���UZ����.��?e|� Ø��j� x.X��zH�k1��t�}�r���|�-�j��0`�k�|��]8�Y..�IE�Q�#���XT^ߙ��f��5p��Q���z���'�{ݦ8
p:d���81��ڰ�,1�UA����k-M�&$@�I�*v�׉���9=�7^��xv��p���&��� 3���׹.vl��~���\R|�T��х�i��NPԪ�\�4�h�N�
Kc�֓Ml��8T��b���4u�����D��]����6���y�`'�mץǎ�\���_,\���&4��j���
%: M+p�"��f����q(fF�w�/X���~�-Ơ_���0�0��O�^�\W�}�͜�{��X�(����D "yg:�q�A1���{�����5��P�����\،�+]�a�5�JE0�Ê�rgw�C݄���VS`�">ua�D?	/ǈs0�jh���#v�f�^��έ�c���}��ݔH��m+b��t��Z\�x��#�)Y�n(2~�t� �RL�H�Ƕ'g�f���O�!�H�m;@ԍ=z&�8�Hw[1�?:��	��0��[�����qS@��!�P�,M��Pl	IIh��D�y�#��|���i�-�y&|O���0���x�k�3V
ݑ닻�w�F��/?'	�5��h���pe.��0��!9)�����4@�rNy���7{����Ka���04R��I2�z�t���Q�&l��4db��B5���Ġ7��u�Ҳ|�ΧeĖ��#{��{ێ�W��>�uס$�4����lC�vx�
?� {!��9�\|{�
�d�C�%���#��l��[1�p̨�ݦ-�qt:������w.�F�����}@\�)oU��<5��J#�FG˸�9���˅Np��	x�41��%{=)��+��6��,�!�']����ϙb��=r\�[���%��v�����L��q�<����*�T�����?<�� ���9�|�
��a����0�T�J��KS���f� �+��� �n-�-� 7A&���fk�%C�-�2�!����+�ipc��mҝ+*I��g덨���>b3[��c�a�i�WI�=A@7nFe��S�����lh~�cZ�FN�������=A5��ֈ���s�ߙuOc)�i�c�x��Re�et�=�w~aȼ'�}x�J��4�$����yf;6ew�
7z�(zJu�i���e)� �dqTuD�*e
�r��vCVa�J��}ʺ�����3W�����L\�}O��z�!胲��2bA�B�/����+�0�h'W����H�=����)!�ʊR}���;��H�`����i�V[!l�� ��STi%"э�ʡ@�6��I��2'��l�bVg2�}��%?u��]��:�Q����Wo�[�F�.`]�
lYMvս&�/,��,<d��}X´��_Z�X3�o�Qi7�"K�Y#���8�����R�-'�$,�K��.߶�7��\Ϝ�ډx�V�����+�z�xߏ�,x�O�Ypt�ԩ;�B� kK(�.vx��n+�P�2��9�1�B���q3�}4��dCѽh68�\wul�+�Md��v�l�hB�Svx��{*��?et 5)'6�_�p�#��ywI���p��~
 w]ũjeI�(�XA�(��{��F�jX��՛hTA���h�r�Sp+!�A��{�����(�ن�+V#�
��{��&�b%��|=,�;pG�c0��_��o�/&�uC��[���A�>�,�K�!�.��:K�m�L(�]çX��	@+R��@%���]Ï����Y�PEu�/=!̳@�T�����`}Q<U�8K��j����r������������0��;غ���?~�t�墺AhS1i]>���8���H����z+:�Zv (ԃ?�9}f�t�r��T`;@�{-t�zc�q��{��Y��Ьbb�$��ǐe�R��~�
��'1��E^����Sx=cW���v��?���*�̾�p]_���e�B��~g�������z��*�Yx�W�v�@�M��\�8�L]!��|G�[�J�3Xۗ�a��kޙ��3;+�1qf�,�6��aQ��	�0��ְx��Y�X^��D�F&����F���H�NǙ�9�O����&s����f�D���~�W���ा�9�cU4]m|$���t��k����.�%υ���
pV7�6T�g�a\��](}P�D�y�k�-�7ߓ�h��P�z�tiwu�$oU!%�/�QO�H�ܹ�"2.� 8��A�Q*�N��NAfK��G�[�M��0���p3�=8}���q�c���F �>�����׬>Fc4�YV��h��z��D%g3D;l`E ��߉\.�6�ĺ���;�Uq�z�@*,�B���AO&ZH?��_�� �ӿ��������u�wϲ1�E����Qa�A��f3�xjW�﫢�Y���~8�g��b����ux[�]w�����I5���t_��(�#|�p�B��=�8��^���0��g���=0�-d���_᠏o�c"]�x�T���Q���Y�	b*�j�x\����v8��C��Wr�ʩ�ל�(*�ɕ_7���nTc��2_熦���3E�!˩�E��v6G�~����-�T���?�Ʀ�*�"��������'	ǎt��M,Р!� 2�0=k�og0��[�Ikϥ{��\��d�o��Y7��D��}>�r�Ke �Zt�M��J�w�j��s8%���s:�v�N�q2���9ӎ.���.H�%HB����-{Kdt��(��I���ZV@UMcs:�İ#ߡ��V�	�=Y�Z�&7桀�ڵ�'��"�U�B�h���O������j��Ku��x��6]�;G (��KS�7��X&�gQkVl�=�1�x:��!�q�o�Q�K��+��!�d��+KX��~����}�r�{e�ន��ø�V�^��n����vPG"u��Ť8W�j&Y9�HA�y���*��^�������R�nD�oW]���38T� �]�;ȃ�,ĂNŞ8N:�-����z~���K�bqQw}P�ĨU�6�E�x�%���8)���O$��B�O"��#a\B�W6�tm�4a�s�b}N䲲I��n�5-W\�M�jpe���T��S��կ�=���Y�� �o�/x��/�lQ[�Vγ��m ��5�����J��[ԂL�lc��")��@u}f�Z=*�r�;�&���/�g��P6�L����jBVG<�Q�ti8/��v>���۪-��T���z���aY� _֞�n>�(���+�
�ƚ�B�:���x��Ii`��gV'�Z���yEyڿց�ۧ���v��,����Q�g���(��o��uc$�l����j5�$Ő�H/"[��"�Q�!-J}�1���)3T@sL�+'�ؕh���CY��Q��y�����ݕ�hJK2�2�t��qɨ{��A!q��]^�s�i�fP6�����8��-���fg}?�V"�d�
;�b2	�G=Pk�c��G�p��@Wml-�Vi�X����]�@�X���� ghՑ��rB֝�2��
�_�*������l\ů����9�]ۯ̌DF7v_&R�����$���DI�t���)�+9�(B6-��ӂ{��V0Bſe��/>4�#yB�rEh"��w������C.�1�C�R�����źb'-nj<�H�}>��B�}|�7EE���0)�w�Y�׵S3I@;�f i��h6�svJ0���
���7�%m5���'��J�o�]I�X��f|����2ޓ�f�N��8Y�>ў�,f���m����(MRJ�o_�:��x����=*2�Gj�F��bpe_�k�8������ �����K�#�a7�Zn����i� ��̹�ߟ����U[Ob���K?�v����^�XZ,������Rw����8N�}��ND�m�t9�4�u�}yb�O�3�ҐԬ����p~�BE���Ag���.��ӭ(�.���Hʻ��<;�z����R3ev�O���)cZ�@!���8AQ.r�m�ݧ�2���c�*+@V3��_Z.\����7����ݥ�/��u�R���$�G �����q��g~ú��)��#�[�5dH��RRc@�l�77��٬�-,Kר�qGv}��@�_�۟p�^Y>[4�8�qV�/,�J�V!P,h@�%��y��.�z&T9R3!����]uyUD�
���h*k�0�[�;1��,Q]ێǎ7����u�LhT��B�DH����k�͵�!TC�f���w�0P��vq{Ss�����!"o�v�,�0k�$d�.� ��x�`�Ȼ��ָ�5
:1[1����,���2��"q	��m�Я�Z�K~� k�s�o����=Q!t��Ҋ�
=� ��C�_'�K(Ɣ;X����%������p���B���貴 ��� �^�����9�s�a@�������.��ڂ��N�RJT#�a�|����e��"s�l�Gv���"_6�3�Y�IX�����@ P_ͤv��q����T���|�2�Q�u_8MW�J|����&�+S��VP���*���Az"��GSP�KUpd�!]�3�� ��[��J��f�bo˫�o�w�=��Յ��St�0�?}I�s)�\��|��q9uT�#Mv2w����O}��7����B�Z�e�6l	��*C�G��}�ѵQ����0D����������y�2�����?��ú�<U��^�� ��V����{?	wDr���
P������t���E���
�0ԭ���']�%�m�<!|��?[-י���\�`�B@=]Ւ�A7�(nI��@L��c�P��x��B�������xt9b�`��J�W��6���	a�����x�4٩�����j�$����]������\��O�t!����wS0�|(�B�d!���[�������>��c�G��9��c�R@�JȲC��>6�W�x#�S���?��חu^�.5�v���ࣗ��M_��$Ԏ�v�|!5dg
�;QU��N�U�2!EǪ�@~EL��Q�撂���K�GY����l*R�WMg���R�t�7�&��y�7�
ś�Q;�f�*�@ᮅՂ`�g��1+j4�I��`���A܋y�:�Ѡ��F�.���ܣA{-�Bh����d
+�{�f~
�7�kf�C�l�<&�9����Ժ�	�b�d]S�#͂�	�ޤk�
���:kU�����RQ���y�F���UtQ�� ���Gs�'��-��f�>02X9��Nn��年2M>KG�oi��>��{Z�5Z��q�Q!�*�	�,�R/Cl��C��(�:�8_����z�1��-1�Y7
&�D��{����|)[�{�f�����T�~�pX0�dQ�� _��$�[���X����hF���H�Wѳ��U7�L]���I��)I7�\Wi@hA��O�ҙ��J$���M���Zr�Dma�@�Y�3Mt�ն-�k���T"xgP�2��^��zf��]m4��˗{�3;'j ;�l��kv���=[i��WM\�P�+��=��Iw;�:Y�ٸR�-��ff �2.��]）Tda�n�Qi�� ?�l�L�F����7�O8�"�p�O6	��d&� ݇�:���ˣ��h-�]H�B��13Q�f�+���u�bС�F5z��WNG<p2��]�ˋ1��D�l;�h���2���ץ�PQ����ȸA��$;D[{~�ە���v1�2��7D�sP�O�K�����ǤIKv�5A��^�Z�$��uN�"Pm��H[N���+��|�xƩ9���N�Z�v�J.8?.�Qr�'v�l���͌�4��x�A�m��Tk���O/���K|�����.��2�A�-z=��$V,W��
ٓ^��:XJhZ��i
����a�_�幐�_aK���3�&��������O�ށ_�K�qڥ^׏-89�W� y3�qo�FH��Bd��/B���TZ'i$5Ѓ�mT�
����9��uiip�M/;{��4��ʤ�Hj|�[Y���(,-�vs2���Lt}O�@(s�I�H���vw9m�[��ڼ�ծ$&��Cx,��3J�R��4�;�JP�I����m����!p��#RU��b�<K�g&��78Eм�p�oi@'��l���/���B(�LyI�
�	%0T�^p�������O�T[�=R"P���u1�ny��s��y)feM�9uT��mV�P	T5�2?c�q���Zx1���7Suw/�Ƹ���?�|����T'DwG+Ӥ���W�H�%G��I���-���|��B
k%.g\E���w��J��rdf�HU%J����_��.�\nԂN��L�����be��m�6��.L�lV�F/�����jHMe_Ӈ�R��ʡy���>O<[P`��Avo����|�C�x�Nn��?c�
K�2�Г�Sb�qH/
R4�5��H�_9w�7#����\@�N۶�{�ƾ=�M4BS���ֳ7�R�yw՜�j���1d&B&
$��+h���P� {o�+ٌ	ǋ��