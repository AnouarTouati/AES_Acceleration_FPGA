��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&Ű��=�b��vT6�4��fWg)l]��@��7�B݂Dۉ�{��m"�?N�vod"��Yd��3�=�X��"�(�1ΌbjSp����"���`�M;��ZP~��B�����r�<d�Ƶ��M�%��>7o�H�(@��ߙ@�
�̠�H���1�Y	 ~����W{��QyG���*�3$�5'xX�}j}����C��@��U]���^�zfgɦ��fA\)Ə@������|7� ��9���J���H�PrG+����皵?{��8�+4�gv��Df�%b��)�K�PQ�$Zi�D.��r1��Ta��M��.`�7 "�6����^陹J�N��HI�RS����[�(.���nHo�s(=��$���n�⺮"�X�Ǻ$�J��H�$������aq-�����ƨ4L�*W�6�V�r�j��6Gv�E�ѫ�����\�x��\�d���h��J����%^ȏ�����?
s��am���N���������y���&ھ�(��0���;B���y��x��r[�e )��NK�9�]� @Au�+Y0`��p�Ry�,�'��	�B����1�1�6,�)�����OȠ���'{�r
��Q]4�J�
����ŉJئ<�VC��0L��9�R�x�,�Y���%)�w&�f1���F93��_b�s�@@���� �7�#=��ܰ�\Q#�?ٚW�w�x�. Yad�,*�����i/��>�Ź�H�~Ѓ���͕|�8*'�hT�̼b�<k���]�C�ף�L�6��[	�X*����3Jٯ�o���_Do��c3���! �$:�J�}�&-��/yʃ�VrG)����9g	
3�}p�(鬁賗n@��|��t.�+�c(�V�݄;ĵ��_���&n����Cb����ߓ�k�Q_��;�q�u=��e�L{es{�R���Y#��Q�����d\I�
�j�w���8�� ���)�T���Q}�U���?\���kU�&�m�^�׆�Z�4
���3�E?�_�_�'�����ȶk���0�C~�eI�ˠ�B��5�H�>��۲�/��:��y\���j�����t��(���|x6�!��Ɉ�������k���M�D�I�AjE��_�ɌG�r�ͭ����S3�7o������ 'ο,�W?��?6|g�	'!H��z�/n~&�8 ��,bK@)�^�w��*�����;�19���_��1~:{��a&:�F3��k�ˡ�V}F;���4���P�`���c8����Ř�ᱦ`j���+a��U��RRa�l
N[������չ:�<�M�l��6������ޝ�a����1��&4G#��=�\���W����O���h�Q˝$��!T�0�Z^���ת:"��*j-=9#n�!B%�.�eO=Qd�y	i��v����
�r�f�j�by�4_�v�#/l�\���]fL�!s�(���>6���G����&����e��ٹ��E���B��o��R�r����i���J'݊3Ѩܾ�ˣ�`����_A�Dm��0F�jУ:�������H�{�69��f��\�[SIa�9B��\S)-�s>Ą1I����y�
��6S�}�+�g�g�(�e�H���} 	@�E�ڣH�(���a��]�*�},��%���qb�6�0�\�k��h�^lE�ʔ�Zn�=��w�� �c��<'i�؟��E�Ͽ�!H�����כ����l�
�'�b}�;�j�Ƃa7��Ě�c�X4.w6.$�L"��z���^t�`6�WK��F��F���!�@TA^V�\�.��W̟�Pw�9y�G���R�P�B�C[\��O���+A�V���l��֩)��GԮ��O� ~&=��U��Y��S����M;o�l��z�4�ʗ��T�wiw��o�i�t�<*���V!�դ�ϋ5a��߅"�y�꾧�:����6GܤT��շ�݀��2�\�Q����@��o�א�tS�����?·H ��4�3�Q?�?^M�-n��p�����ɝ})�����#�6�VA�8�\���[&�����TS2{O�b��^��PRX��l��md��_�d�Y�'���L����M3)�O�z1��m%AU)�L
� �+D�:�f�4����1�TEw�\a>/qX����=�~�ч��@�Y�#�o�̄�V�CD=�s�ha+����띊-F��қ��'���+��]��6.�a���x�V����n�X���`��9��V��?�!����0�ėqT�3w�`gX	<l��-�'�o�%��&��G�X��Y}�DyUp"�k�	èpfÔ�Z�}�Zh�۴����z�f�}e��A�y�)�#�}�;���Me�Ǖa�kG<�L��H�u��W�zrh�,swq���:g>��֣���<2���&��/�a��3�R����P0� ��l]v�BcwSL�%!`�ؓ�z]l �$	��ٮ��69Ʀ�zqT@eE����s��V����t}?R[�T$�掹��jٺ3�L*�͢�A��9��H z��*�4�� �p��pP.�D!��/�H>�5�
�X��=��3e}��N�Hm��f��,��A2bX�s��g��(l�#�~K��!� �P��`�31/�u�7Z^���:�7�m��e��m)�6��!u�~W'�U�n, 0Yx7���s�O@��R�/�I���I=�M;��O�[v�Y��?��t�������y?��3l̍~F�2ܕ)HqeK�02�*��6��kC�b� F�1���)k(鿮f���7+�\AѬgҴR�I|�:A��ذ��S>��^��_�k�?cUv�9<q�:�62������D�7,B�
=�qL~g��G' �Dz��kEc,��R�@��7tt�;��I#��
�m���/x�EL��N�ߞ_����ѓT�*���i�I��+�����Ș���y�ո^�<{��E~�مV!Rv.Ye�]5���H��yT��`����Q��g�i���?�)�,�.�Ì�������$��c_���Q̎���L��p1_��|�fm��r1������k����EL�F���������P��+�����Wϼ���(��y��Ȳ�F�_9���I�J���2Bx����n��fkN�ʃ�v �7�I:���ݹU܆:s��g �P�2��E�cSA��L��@}ow�����*�'������d_��܌ܖo�=��DU	O�FI��yA�����g�2>m�L=}$��7�)9�&����^&7�pt(z^�#�j�Qk��̵������;�\�D�1K)���y�� �Xn	��g���������z:%s�/�����|d�����p����w��M: 8�}M��h�iG�X�<^�-�Jt��HNJ�U5s��q�cU�C�B���0S����P�e���*u����=�Se�FK`5�A���Jd�_���������P\b:���5��R+���M����ȗ�/��� �����C���G8V��Ձ�8��p>�\�����dWڼ-q^j�|As� ʿJ�m�)��r{'Ԓ&Z��G�͚a���P<�!3[��c���10�ب@�O���Rs8TP%Ss��_7�0�i?�a*kR�m�Yj#�E�A5���o?�/:>�b��4�u�
&'�A8��`Z,jψ=_�"D�k(�`)b��'<#;�Z��g�Q���6I�|c8���<6�\�Q�M�XҮL^OP*OFh��la	 �z�ƛZ��4Q{e���$Q*u���o����F��:��X�׶�4'Gy��ʓ�Ӌl���X�	Kbj������+N>d����:�J>�ZA۴�cQEjk�f��j�~�3�Z�<��f����X�Y햏�L�u2Ә�ǲP�'��q��Ƚ;�n�Zը�Ƕ&N�S����b�+�'�{B����M��,�3��:u��1ު��Ӧ�Ϟ,����a(kr�v ?�)|f�ޏ�k)`.w�r��q��~���Y��d+�����M�ҳȸ\��<��3�����>_��FQF�%:�?n4���J��xE�&Bu��r�d����	��_����J��	&�ov.3|���K�{G�y����*�7@��6y�h�
�.�zWۀ��:j:�������&���??�:j�Of���/N�do���t����tACot�ӫ�6:�io!_�hpl1���4zU����Ԕr�#=A��_�}b%mqP��T�O �8
�B�Z�}����B1b�k���o�@�g�_,1^X��ow��DX��E��O�O���;W]~ik�����������1@�O�˶ Y���t�wp�&����=���c�0Tb�h��,5��������3�@�@ ���	"�v��zJ-�%b����Bd��K��%ūsAV�� �3�m�g�<������2w�E�_�y%�m��d7�?-��x0u��KpJ�� ��T�ʽj���������\M`�^%8"T|�s�;ǴD�� 4�JU���ڈ~��H?�	�S�1�����W��Xu�Y�E�z  P�B���n��K?1�8��m
�END�$"ϯ���ڀ�/�:�9�N��ڟxbi�Z�ph�T���^(����-���!��آ!;��w���<\1�*�8eH��|_�ZDջ:O���5�@/�M�I���/}x�.���z�䝭���@�7Io�8�)Uv94=~�@�I������{��yTN2v[o�G8"�&�?cS����1�u����ܕ��@ w��S�\;̲
"�s�9��֞����lT�7�|0V���r��+�i:a�eo��E
[_A������I����;���;^�G�=����m�aԱu/<X��7	`friZ�@;@)#]�K�)?��A�~V^j�k9�8�?cc����X>�?�%i��®!��p,Τ"\��%d-ȊT�fn��;.�Z�s�#��Y)�3�O��e��-��b�g���G���ё�WQd��tR���4^����x��Z:!��I��!l�0V����1�e�Z��/�ˣB�V�5��8¨}N�O�$�B��N�*�
��G$dIt�w�Vl��d>I]����b#
��)i�^7r��⠟�.j��g�*kvS�f��#W^�3/>�,
sN8h�j�F�1SX���m,��T��V����$�K�J�%�@�fd��Z��Tc��Ĺf7E�x\p/5{C���|�v��`n�N�I2��\K�D��;�k��(Ođ�f��ot	w>�tk�����Ҹ�9�b0�㋣�e*v�^���C�8�~o��/P!�M[J+�fȦZ�}U�X�z ������Q;&&�x���'���F���Ԝl Q�j�s���zC �~?�)e����N���I�ҝ����f�9I��dzB���ccvw��+۹��iL��0:��6�hw�?W7�9���W�z�H�>�&�/ǙG��@��Z'rr�ab�����Z�W�q ��	���� �>�����Qa�F5��ы�����_��&ߴ���*�����I�m'�d�����D����lTh/X�: s��H�Aa�)�>��&�6�K��Mb[6��q�7�����O��`�-Χ��c��y.(����=rA���(�Am���VG�bC)�h6:�&����Eo�nތ�f��
�X����$aO���L������Q;��f��c��*����3L��c�G#=��&����T�q��d�?q .:��3\�&^H>I��{� ҋT�~��3o�!d��Cͅ��}�i�&�π�R\��@�ܵ�g
��[�Լ�:�O T�9X�>���_9i��#�?9@�1�h�wg�V��qXMfi�����O���ibHى`�2�W�ͧ�݀�Cp�VU�,S�Ms�x�x��{��(���A�1�bY!��J X����a��u�^�"�^dtƀ`/��̤�6]G{�@�L�_'�M׵sR'z"|��x|("�)a�X#~A[��d��-�yr3tW�'�7-Z���:�|n��T2	buA.c!���6IMP�K�ȨMudt�Ĭt��ː�x�oW�յ4
�!{5��,��G�(����ڮ��+ �j-`����&$۴W��^�����P�0S�)��� ̒��*�O�$��-���H�X{?	ˣ��I�c~Ā��'G�l[ �G�Q�c2���]/��>��u�r�=V��sP~�>z��CV��w�Ї�����ݮ����iiCP+��?�ab�H!�����]J�/9�VX���(o��<�[�T� )cs2s�bIP�cӶu�[a�5����o��JA�E\l���O60�4�U8�Ɠ	't~���P�)�%��r���]s�`6=&��G7M@d�_�C)k�Ws� R���"K�� ���M���bJ�����K�vaΙ87yI$Ɩ������Ң�\�+8J`�����D�8��1;�I�D^w+
����+�p�ڂ���x�]a��Qs�unFT�t��kz���TT��Ԝm��^�8\Z�����}�y*���t��(�Ît��ċ�է>���D���д����&�~�}N��o���_�W�:�ґs�PZ�IX�l�8�d�T(�6Kn'�vc��}�K�z�^��;��DOw�u�֓ D�[j4K��; QŨ6��ba��AY�{��>�3j�Kl�/�L�LD�����V�Z��V�F�DA���yC0m"������H>H�N��4���L�ǰ!�P���]s&рn+�?g-8s��L�j@j��}D&�o��Ki���9[��Fy*�vQC�;�=��vbh\Y;,�w1�O>�e����z�@�R�4U���e��ZD�,3�a���|����}�ɤ_�;`. ��%HX<Ţ,3m�I��JK���_���=H�}�*�T�"&y5���b{��V��CU�)ᦴ�?U?F��?����V�P/�伮����6�q�|��{ޙXkVVϟ>��qo��u=s��'�2���q�\�[nyd E��=vjL����-��p,���k	���mXOCThs�s�����ْ02L"�O���~��z��kﮋ"\SY(��kq*�����I��ӛ4�rEn�	J,�R�$E=�I�+L����`���'�xv�3%����_(,��g޽���&@RU	��D�yݘ$ف �O?F6�ɼΏTX�6 O�@�dڍz-FͲЍ��x���U	�=m�!�6J��^|#Ύ^K/�3_"���.:-ψ��K�/HV��b)'��K��\h޼{-05����xwZ���z���^�������M_�Ɨ�jǁ��
oe6�H�8���5�~N��ּeMG#>��IѾ.�_�Q��q�$O%�CR�$(h�&<�ί��u�܃|����X�[��Mf�L�|�g)A�Rq�l��&�(�O=�����B�b,�6D}�fiwƉ�f-ed�|
�/��P��E�E��ʿ�	�h9�-%g�X	_����Y�����)W>թ��!I��16�?�y�S��kܫ%|0������'2; �{��+.��̉� ��pm3�+|�<C��!��W=��߇���}�)��xw�!��c�e���K�J��FMO�	�]�~?Q���Ft�H�\�ޭ۰|%	o�	���֢��]2��3y}@���/Q�g��7�Hd5yC/b�MVJ�Y��{�
�Ki1=�xLΥB||58�M�g��U �Q8�!�$��H���.�N�[�Ϥ��"~ʤ����|��f��h)$�;.ߌy>z\zK��[���oL���`�g��T��c�&��&�?�{?�.SRf�3���v�1x/r7��p��3a�Œ&�|#��o�S�2��Ub2��g�@(,��I@D�̟���O8K=�� �C�}�?Vvᚈ��n��gA6��чb���
��L��3�ړ�rו/��fNh
s	�&ux�N�T%����Q�Uߴ��(K髕1p-�il�'Z�����L��C�*���8�0e~�3��m��-�����X�0�y��s�$s�k揼=[F'��q��+���^@�������gw�7�>��[B)�ok��G=�@&�s���M�\�OK<��8O�	�\�^�N#	�����hRg��G�`0��B�f����6������; Ҟgz��I����m ���%̻�I����/@�D=m7�غ��W��&��sx�0�K�(6M�6��5�e��f���P�6 �q�닽 #�)���6m�dc��>(wj'�A��J����E�O?:w9?9]$�d���|��^��@:�d_f�-����Dy�(ؗ;&��|(�er��7/�qK�>����n(�/�x�Dl�.ёE����^�/ӒFS_Kq�&i64{�P �_�g��F_��+x[_,a<t1�/�	����"�s]��?SM��VEZBʙv@X\�nBq�����L��KN{�$o	,>X�ڵ������ x���j �dll�
Wr��pp�����t��_�+���>g�]��Tgn!��>9��69� ��Ǡ
�'�� ��Y	���!֪��U�f^�3�} ��ڌ��Q��a\��4x�u%�k��Ab�X��#O�p��Aq���<ϒs�-Bخ
I�Z����59H"�2rL+v�>]�}2��Z'j�1�^�A���9�p�MDm��ɹu�?���p����ڦ����_O'�t&� ��<ss�������ݯ�AG���<nFb[�v��qZT���I����ȋ����N�L!Raϔg_��xWe����'<��B�;��_�:c�L�J8L��1QAIg<w�l{�pԹ%2������z�hY�^��b�4Fk���vA>�'+�S�_X�6B 1��$Hpiޖ�����CZ@�X���?~D(!a��c����]�\�'���+"H�b ��]����S��@�p����F�$V��̅BZ���ȕ��t��O�m{�O���]�.G0� &!l~
-��#��񝞼��CXcPo¤U�=�t�;�-�؞�K����<�rX��\ �����q��q�b�K�N(y�ݣ��<�����'h�6���-M��v�W-��g�9��q�%���MҘ��.�����1��f1�\_�gVݹ��nn�8R�7k��҈g�����^������}^���eܯ-�Z_d���ɜ�i��u��k���Þe�!3��J�д嚅�c�	Eb��j���9`K����lxb��C�N�}M�7+�/S��@�g�+�X��a.xj�zg����bV�xX�3�J��S��񹖓4�F��x�����U Ax��
|ªx��Kk��GvQ_�u�-�H�U^m[F�q�x�1�)�D��ڧ�.�q	�����ݐ��
�7�qI�B�����DI�2�����X�XX��kF���{bn3/�ܩ%s^b=,�#~�����az���ӳ�_��(^�9�6�7����8-1ũr�H��k�?��CE�� �����>�.����/��().���CN##��1��ƃ3 kb�����seN��#?��2g����Y�����:����&������`i��8��7O̧Ŵ��5Ǐx���	�.�U�L�"=��O$[��Hr��@ޣ��m�lŲ��Ɯ��-�?��>�C����ߥ]L�s�Yu_��*��������2y���^���[�&��3�Ho��4`��Qҩ�Q������th׶�k�'g��l�-툥 � �F��@T�x�K	�<d
Z"����r�df���,�@��άҵd�g�-��J,+�R�:xh�>O�.di
G#%��6���K�s�A΢��ea7����S?��%i�n~�1�&���ղ5D�4��$(�_��Aٺ�M0�{ԫ�%!:{@�q��q��Zʷ]9͉�S��T=�B"Uqer��@Hw�P��c�f�ק1���*���ݿ�*�e��ԡ���f<�����`A���U$K�e{?�:��L���>�w���?�z�KT��o͌��^�ɲ��g��T���*#z���hC����W��C�r��.��E4��`-{3 ۝r ������X��}XEW�6�o�#o�1�_i���]��9*�I�\�/"�.�}���۹��a��O�0dMl_�Խ�ٷ4���������)���6P/*@��B8C�#{�+W��F(�^�)���<�'�2
VY�0A{�b�n�8L�d���_�j�*E��si~:1�y�:��{���W��6GA����X!zɽF)nA�Z\�4�]���P3��2<�R����,�ȱS�X^��zx�oP}.`�$Ԟ{��/��Ga��a�ZF���7��m�U��0����{g��F�Ɉ�0����4n�]t��j�;�.t<@����>T�G^<�;�_~����]	@wR��d��qt��h׌��^+E����4����,M}��F���,��^��~�`��Dp��e���v'׻�!+��:�lʗx%�Rjf��M�s�g.����K��v��Z�����G��a�:&�x[����bĒ[K��?J���f���f���W��?�ժ���5�&��H6�]����T��6Bx_�� ̃�}�8�w��	ny���㴥)@XLP�O�Ŕ&��!�Qr�k�i��d�Z(���q�����J�K��C�,��:5��S�3_����8R����a��j�j��Yř}}-�X�@R��bхb��~P�?��O�)�~��g�Q�E@�o���┪[bT�t������Qc|o_�F��Blo���0\c��\�͑
{�]W¸�_LF.���C�T׾y�����.���Lk-B*]m�`�<�,��ӷv��i�Y_�Ee�������7~�9c������[�tˋVO��u�i�<|�t���;�VL����E�X��i2�9g��)ĩ�B�9�~����Z\c2�/�0ၹ!<0���X@�z%�c�/`mH�� ��ea�QW@�I�ť	,�k��n�l0EF���#�L��,K�=����_�LNiI/_��9͙xe�V�yT
�
S���o��M�Ҙ+/?m�{���i�Y�n�0L��s�� E��/ޏ�r���>�Fo���vw<_] &����7�-�}���Bo��V��C6;���O~1(����9�EO�������/�9���ME_�=���h���.b�_�:u/pkU��7�5��;0�^U�E��/����(�~9�>������F����/�:Y1���r@��&Z��8���C@R��؜*w �&ἔ�G��FC!�l�JGu��ߓKs���c��)���X0?Y���x?�Z&��IV��;��]d@����L�k<�b�:�5G�h+1oEmT�$ �;l76��h0�}Z����a�=p2IJ�I����rUa�{1��.jL�/T�o�]����E��E�^?C�9>Р��ܫ^��A��.�q���L�j���J���Ft)������_�zFybc��i��|�Θ�� �ʪ�[�TMhN�����̏�j�Ds�Ȩ����⏸��6������%�b���7�Զ1z��R��(?�s�iAQ���,��
tM/``���U��^�f���f쪤~�l���]ࡿPg�1��2��=a'N�&@-��j#��s�_���{��������-(hM@��QR���3�*�P��U���½��Uy��%d'dW?��7��h����#*�G�C=��ƓW�V�����`�}��i�����K�$�"$�ܖ7n�K��:�����^�-˂��|_𮦨���~c*/��\Y���x�!]���?5�6�1w�����Dk*���9h�\w�;g!]J7!=��Uxh�A�\6�	EB.����o�Z
>*�cf{�ǲ�W� ��1��"�BUϣ�x��9��Q�@,��m��"x�H��u'�%��`��O4ǿ�N$���������H����3�$U���[r�L��K�1Z���בJ "��vIF�_5I�g���ٳ��c��	gA����X3c8�A����i��%�n���X�[�n%[�1�ffN��������Hi�P��Rt2/��L7x=>�__Mw.ۉy}�D`b(,��(LBnuK�Y�^M�Tc<�*7ޠ%���G��?0�uL��wb �{"�V�FnJ ��'��jd3U�(1X��ºg�E�C��9 P��:l��t]�\ �aݳK>V�}��--�?Î�0�r��:�� O���/�5�ty�*8.GxѦ#�ޙ��r�;A���_������ig��Z��)J5DҾ�u����՝����Q�c���?6|�z+��5��� `���o|7��N�l�w	���j9~X�z��|�֧�����b.�7�]#�F��T�q䄴[z�w#e�Oi� �ny~Jw�<a�dQ�*�l�~Y����fN��LY�4g����6�mA��CM���>�P�HiΈBWzN�@�g����df���q���1��-�����:��*��3J�tF>��\��}U+���MR��,��I�v9�߈�F5_��$��w�o�ѺXTl�Q��+W������w=��ױ5��7w���z��D�Ʊ?L���b�H��ȿ����M�4�Y�X:MM{��J�'����
�H�7�@�I��s��jޞvA-%��k<��ԟSʹ��lOn�g�~^j���A��cRt�Fo{��q�ѐ�xK����ͤ��E�~�{�g=��<-�}v�Ҽf���)"�����5<�Z�_�ɀ�e �<�	�����1�m��O|��c�n��k�\;�� Ϗ|}Q�0ɻ�{�Qx�&��� �(BSa↥�uś�a�V��㔛��I�	�r�ʽ���2����w�e-�2۾�h)�	;
!S��)�V1�U��]`�[7�g�iP��S��胡���|Y� wN��:HFD��8Gzfw�X�N�>�y���8'���^�e��\�
q��S�1G�J1��47�0
,D��vĘ3h�D�[��#%��"�j&5�g��~��E�,���4;a�l��e��[�o@<7R���%�:ˑ��G�'B�r�aa���� /@ޅPJ<*M8"��+�I���0H���<��ڏ�4�-��U��u�l����	S4N: ���<W���ǆ�!b��z�sޯc�R�ސ"��O�9����� �Sj,�j2gS�+:�{[ƙjn-����H���˅Ӷk7:��?2Dt�2T�C���'v�~��J�KU���^X��̾��dk0�.t�W��X�ڃ)�	K���-ύ:m(8(Z	K�çf�|�rj���Ϭ��Â=:�+[��/l���ݍ�k,6�F���5)>����=5�JѤ�:;�sY�+c���[�/B�j]�}����٠A����H�����t��s��d�C���ƚd	��Cl7�s7�T�؆���k�M�ݔa��eCp>v>l��aԸ�w�.���FT*�%u`�tf$�[]%Cnge�����J0��r��)����u�Ҿy���n�y����`���A�t��ӯ��R
��<����]��^�,.�k��@ge�%"�Z�A)����0Z]GW �F�ԟo�K[7�F(��~�����ȃҷ�+��#37q]�!\���u  �����b�`���G_��+����˱��B���/�+�9��^g(q@t����>y�*M���>��}�u�"���D���VF�ڷ�|�t��˾�{�O�.�F.�YGV5�UN��q�VÉ���*��V�(�C����%�re��"<��ظW�0��Ç��n��s!��aP�F������-i��,��O:}s�UrZ`a�5��:����e;H�;���W+�MF���4�ѕF^������R4*&mE��]$�w��F�S�X���*���٤׆�R��,��46^1�^g��wL���e�#<U�c[���$G�2�ph�X�K������+�E�Q���Ϯli�]T6�a��\�G!��:A �# r]���}&[�Q#)0Ce�<���ءM�^���O��Ͼ�&P�ޯ���t�E0�X77~�݋8�ӿV�3mk� �,�6�'y�#�g��NCյ�h�K|3�1�X���{ٟh���Tn��\'u��ڳ��0��'���@%�^Z�����/��B��皆����j���rL`=&'6�rX��d̳���v��LNޠ����/z�d3X��x ����*#�:6��%ô�������W���^N�x��!=�s^^���-gJy3�P�x >�W�d �t�(1���c����^<�dC)[�f�y)��{��R��n9�Ge����5bg�[�4Cu�(���� #a!��1��"��%����%����ݲ{z\㕌��U1
]��j��М����ӹ�/x0�S�.]Ƅ�Y�(]�E���ς�є�?'�L��Cx��TDR]������=H{>������h)=��M������
S:�㷟��C��.k���x�1�Y� �U�FM��>��"+�LP�"oC�c@U:�c!�}�|��;��0��&w�DV���y/�m[)V��`�^����ɗKS������.�e�s��d1?��,*Ȗ���u,��H��2�뀷�8{ϣ1`Λ۩�A�_@��!�/���"y�E���a���I��f�@��(ʃk�U��	���V-Z�Ș�vp�zH�B��\���d)02���A�z�b���`��h�#͡Ad]̋+!^��ɚR��Ew+D�dm�[�=��U2���V�9Nrq����B[Q� E4�2A�NZ�&�;9U�U+c�����^� R�l���n�?v�;k(F�Cw��m���^�r)�}�q�)�]���~�P(D�"/ R��y�7K�5E/�j� ���0����g+�"ح|;u>�Yi��(��@���|?Sw�'�1�>^���(/���Ki�6 ǳ�5���`��1�̳Ѱ�	�e
��I�d�ƹFb���.x_�6�A73 �j�<9 )��I?eB��A%��B��U~Gѿ�~��@%�M���U��uw������B�\�.C�G��3�yݩ�$���Sl]v�њr�y:�ۙ��:��&��f�>ް߰ ���|��q+jH6�I�	�ۊ�h�"DW��~�k���CKݛ�ky>�c0�q5���B6Х�^-H�_�b�2wO����q�5=r�0��y����(F+�l��i�Y�4}{Jp��a���a[b�Jr��w=N�BOK���Am#��5+?��KV�`��{��o>" �tu��y���ke[�f!�z*Ü}8���Cc��B`1����vw�@�����FP	I-'� 2?�;����R��O{v�Da�������{�\�7��\�V��<����_C�f�(əp�cYnS�Ҩ��e�]4��
�g RB� .������[��I��_�b!̄~�gv��S~���P`�Hh�KC�0z����)�	�C�%Fn,��=K,*��V$�)�0��p���ߨ��6|ە,�4_D�XO�nH
%������閗1���C�rq(�߃���Li5�`a��J��5M>�盭���=@b�ZZ7pJ�$/�#����8�;�-"6�#<�imZi_4�9қ�QtK�C�];E�GQ�g�uFz�Pf�a+1U
���� 醩�#g$oU�b\���)��ل�j��uF��$���sݛh��O}'Cr��H���>�F�2������a��)��md�y�tS��r�D��)�7�I?z������!fۿ�?h����NB�Ծ�+vHr�/YU���Q�y{#\8i��0Z���A�0�!��5�*d������#n�n�X� ���E�4ޮ�Pm�D�-��˺0�`"�8���ϙ���q	0�g��'��Q���s
������yq-�+���V�a[c�H2��}��.��8,�CrVd��c�"���Y"�'WB�l�Ĉ�߀43��ǧa�Q�j��8�M�����['�re6J])����H�2&uCa0	n�x֙LA�W׭+��6��E�H�M�6�<\x�C�k��_������C��Ҙ�b5�u����H��=�v=��u1����R�(/��-����y;�4ܛ3��00b���yXHf�`�-\uﴥ;I���mӿAz��%����}�7�a����שsto@��Rx��M�즯�����|_�F��?����!9���`�)qIwV�ϸ3rO��]���Ě�ߺ��Ѯ/��<s>.d�"�h�ۻ��*���!��[��6=��T�0#y�֥4�`�>U�!���=��uϗ���>J���a�Z�3�:�����΃�j/|<X��r�{�.S� jL�6���W.0��R|��6������x	�����'�Lq��	:N��:�=�|0C�Qt��!�Xt\[�EB䯳4��`�3�Au�*$)sP�<��j�����U�	B噥�Lq��?�V���U�i��~��mR�[�R��a��J�!;��v x몆���l��$Ʋ�|:O=o�(�Wev��(��q�Í���oz�����
�7�IJ"}�ê�e]������H�b}���!�HK����8@��������|��v��T�SF[c}��� ͼsE"���� ���ōKx6T(tl��?
�����sgTZJ=��S�zaǒO:l��ϝ��)�j��w�I|(��D?���/�4�g�������V���e
�'�,���6��7�2[�������j�ba���u|��zغ�>���ܸ����
�_���7ԡN��b?«++�d�����[�3��޲�˹?��j��T&~Hݘf�F V����G`�IWn�!��ɰR�*
T<?������O
�z��#���,R�rP<C#�7G�P�e���;ّD�����ttv E{��+�q{P]#��Q������:a/�r�)(9����$U�Mf(�WxQ�ȭ�ȭh?{��R��hçm�pb���w*7l���"�\Ca�=�/=�	���A,�����)�I�����	~q�~�jI@�u�=x�:`���nh�3hGY��x���L�A̜�}��Q�l�b�r��@�v���S�T�a��	?ǩ���n;��j���t1��v�zZ�aQ����O��,� ��>�p����j#.�a��Y�KB�������k���Ko�y)~��EN���X4'��r����Ч�#'���Ϡ��� ���4�B4��]	�`�b��y��c���Qi�U�\?ܹ��V��1{�z@��o��Ұ��L8��������dB�c�5�|�s���|�'�{���M�m���q�҉���
�~w�< �ζg�[��[\Cl�Z�����hsy�dR1EE��:��ڔ��$%���*�A>u˅���BFoc��]#3|�ъL�!�k}�O�S��y3�5�b'�:��ʕKxY�I�>�vW���+)51��ב{�>�z�S��4~2�B㯜N�|��J��TD#��_$�F�������l�W^�����5,^�� ��d�Td��~�w�iU2�й��'�eȆ	v���+
z)`:����t�9|��&�·1�
\#'���dg2��㢧�X�S �l���>C�J�߰Z�/�S�Ȗ��8�A��Y�	��@�a��!G(�R�����T�@gR�)�;W�M,]�ck(w���mvҫ�,�E�SDlkOef��}T����
���ґ�y#�ӲAjo���#�ӧK� �����a	���3���_����99�i�歃 }�_��@8���;8��FǄO�2,h4��*(����U��+8�q�/��-�`��!⮈�g�g���I������v"�%�k���N������2�.X�S�5B��V�Z��g �Uwy�@:��}���H/�S<��
!�S�%�P++W}Q��͗�/��H�ÆH�܍�ՆQn�C"��t��hfti�n�(w�$|�&?��ԅ���yr�s��	Ա�ՔB���˛,?˜teLA��>c:~r�|���<~����_*��%W;�S�z�$d8�dCHt40�oK(C�;�-�;����>��t��`H�a���(�!�W>��ޏ��O�kU�h�b������
��� �Q74d�[��cId��
\�W���նǷ��l?F� ��Xo��K�"Ar��L+�kZ�`�&o���V�W:�F[Ԩ5��{��bO���	�z��X�y��i�%90"d'��0)o�C|�/���	���w�T�2Ȥ�����2����d����2�������fK�n+7r�+/g)�c���\�g��ES柙A�V|9�	ӈ�u�v>Wk�zb�	��o	L-5ese�p��	��Iv��"31���V��o�p``ό@�j�V�>|��7'E�"�y*�5��?Chx�UM7��2q(A�[��Z@��
k�p���&c�b���]	Ԑ����R��dۃpԼ��^��U�Ȣ1�w��1��Lי���h��bZUÏ�rڼg�v����Ǖ�`qE v%�+}�\V���дx�]F]~�"�_�Q���qh.���لюj����}�8k+W>�=e�-<��̰B.��"��҉���3;�A$(�-�l��2|��D|�o�0:��Y������@dW��@)CĮ.Do?i�����7�?nx�2�<NFYQ 2�0Ez �k3�?|K�>��N��^j&4��s��2l�u��_�.Fȝ��_�V>�k�G�9�Uǈ�{�e�kƟs�E��|���/����x��}�ɷ�B!�eex\_{9+[��J������V��]�"K��Ϡ�Bi�a����qtT԰��%2���P�sO�k�����.m�b�R�v�b�4��}�_?�T�P�9"?�/�2_w��4ܚ'S�a;c7��\0�1�X�A��5Y�:+�3d\2_�qD�w<��\�_�E�F_;�JcH��l��C8�`(�o�^!�oY���$u�4�4/(��䵅8$\�0�� ����~(����*��"�^m�)C}I-e[W�P�.~x�4 ���u[��߮���O�)S(Ƀ�IM(�%��^uLNg̫���^����|[Ib���Е��d�OD�S�O�e�#��rX�ޒ����9�w��_qnO��p\��߄�Pj���D��K
n������&nJ�3g&��L�e���8H�����A����hkV׾Ǣ�$I`;(c��R��TN�)lԀI�%��Q4ז��o�3ߺ��>��4j����*���ۉ���kj���;0�4�����$gI�k�l���Y��!V��#jh#��`�H�H���4��?��~��;"3���~]��w|?��2A�;O#3V��A>��N30�{�Q�a��`
�ڢ�n$e�:��O����A�[�1hF�&[ɪq��>2J�m�(�e?Nrg��t�����?h���$�ɐ=�/,���Y��J�K>A�I���-�2�wi-�����N� �}�F{"l��Z]�{�V��3��HY7ڼ��:��K�d�[Zy^(ڎO���~�Bu�"ao���.EZ�.��ڥ���B7&�m�;��8�W��fw�H�2u4�N��ٰ�&9�'��t���)y���猝�9��cT�6 jP�P��a�d�q�¼�8ݥ��Գ(흱�.��Ҡ$��� ����T�z��S>���(��^oN9@sW�u���+L�Mc�����𴙧9��Γ����w��~���A�_�c���V��v+Et{*,*��aXS���P�3ȇ��pV�,B����u�#���P��D1ϰ��r���@HE�[�)J0
䐩;
��k؉d,��Q���uf&�#rQ��E���6��X���Ŗqfd�Ц�P�p�D-�<�EX���͜��oz�M�/�X�ݬ �J���dt�s�qUac���Q�y�_}�1Y��<jNW%��Z�ֶN�|��2�>r���õ �t�J��Q����#�\��@��4gX���ܿ$��M�Ɍ�F� 5��f��&�$}�1�fd
²~����Gf6�%�}@#>�T#>�(^����h�@�.�ҟ���s��3�	�<�&�˵�1'TU�Y��óCҡ��4A�M� ^��/�A;ԅ�,�M��,��w8*�/ߓ4@2�57Hs�$�ҭΖ��dћr/L��4�F��s��F+�_r�c��QJ>�k��h�HP�8���K�=�N-)p��MN���ނ�\��%�*k�e-���{oyqg�*&g���b�,/ZlՋ�����r�����Sq�����\�Z.�آ�V�l�!�yA¶�*�UQΊ��l�D�C��������r�V�S�PI�#<�|k�A:�<�֘�4�#��E*�[��5�Q�6k�-�P�C~[i9u���`�ۤ ��K�o�$� �%��sQ��g�gg��(x�s�t�um�X`	^K*���8��<�W�t��G��^�O$�<K���֤{@~��o+J\����Ϊ��|��e Pw�׮w.E�@vA>�Cb��s�	:�x��U�ǃ$��L� ���y:&3D�5;	�����W(�SM�y8����R��M�+��$5G�q�#�N���' ܬ�[!(ң�>]�ʾm�Y�"s�cO��vo:�&���	�5_z(a�3Y��F%��8Mg��_�2����%��@�[��`J�S��)�1;I�]"UM-�b���ե�f���c
��>;�>�Vn�w۝#5PxjIǐ���RŊZY��(O�F�k���o�
|����?��a���������K���4�����+�p �jJ�T�ucUP-�$���7�NL�[�h�<�8��Pv�/�[�s�<�`J�~�X��!��!�ҍҳ���<R�-e/���üLU�v�q  ��d�3)m�f��DB�m]x�L&�O���੄���4L�D���
'Xm�9
����Wؒ�?���K�v~۰�E�g����+������ؔԹ�r�/Z1,}�S�����1j�0]�yv;u��7�}��[]!��-�;)Bn���p�m��mc�M�$wJ���K٫��oR��Α���<���.��4u%��S9���}X��cc~F��A������7Xdش�)`�i�ι��ޗ�Uh.��R� ������:L� �h�⡸���t]k�}'b�1k;��NN�|$s9���g]04�XW25X�n�N_ĉ�fO
��\�fY
]��d�X���w��L-
��q��\��w|�����7-�:�+̑��F	E��%6����`����Z(hE�H^�=~^��U�+�]`T,��_4e��1(}W�pZ�)*_��}�/ZsJk˘O#3�8�k�jI{D��p��P�AuS[j&� ��pdp�7��#�Z�ܩ�`�202k �� y�k\�`�|0i�����i� �wJQ�|'�Ŝ�(��<������ot������s~zE�\��u��3�����x���%0��cL�0��Ŋ�DT���LK1,������W9�rsD��D��-��ߍ�l:]��R^���)>��Lgֲ�"h=Z��ْ�;g�IE���13��X�t�pX{���� :{Em�\�^R�c>Z�5��B�W)�ΜӦ��-�{�<����.���M�U}ߣ�i��]��5�����D��;Lbmi�������1�qN��c!��x٣R=˟�X��x�|�w��OQ��S-�2S25�#Ì¸��&��¯�f`=���F�d#r�}�ҽ"Q �=tS����PwgU 5�fƮ��w2G:a�63�>o�j����\�_�ꥒ�����z�������¾M����T�1}��+�?���H>��_B��ߌ�b/O]� n�م�hV�T�\G���QMѹ��x�,�ĄO����'���!m��'�M�'؊�]���~N��y�A)~��� B��)!�U D��K	�Y�h�cH^�E߷�
o��Hr'8�L��^���"��3c�2�C��V�3���2�U���	a6�@��ō�X�ցy�X�օ���M��D�I`zbA����ϻ�=r�d��N�ݩb;`7�x�<���EYx&u�Ƨ �z��X�yy_-���3��\��К�$��FT�s�'i�Ȁ4����_�;��e�@z,�����P1���a���|��҅�����Y.�9�܋�«�d
sAQa�T��Q����5z������S��K��b	2�2�$��y٨�T�YƑ</bVfR�ġ:��� y��|��	���{���(<���z�����AJFm��S���KN�ͷ"�8s�Rz>\�Ȳ���C��Q�qy�hG�d��R�w�s����}z��Q�?=0�>�m��6W�Z���>V8{.I�۳�S�;�T�O��e'Y���z�ꭥ#��r������j�
ש���6��g�A���L=X�F��	��j*����ϛ��#1�8�M�u
+;	׫�̓_N|/A0�_�whLR��(c�n�!Aۗ3�0����E�s���Р6�O��D���G�,��Rjޖh����VA��������v��k�4?gMh��]�N�T�VI..��K��˖x��{��_��^xp��\`��R��.�؈��U��}Fp�td*FW�}=L�U5�2��S�����L��x���	�WW��
���;��牸�ӣ��QG���4����}���nU�l�^f���4g�����f"��|n}O�H�f֮3�h�4�5t�nF?&�4��l;����t�x�WU�6�`fW�W�T�Ƨ2� Wo�o$�|����=}o>�Z;�8���K�W�M0P�m]�k.����G�'�������Y͉
� ����.�ʁ���nY�7@[!��g�P��-	O�+K�ڌ�1�p����X��=Nw�&��ӳ�>$��tV�U��欦A!�S���wt}e�ک@%`��4!�#�P�>p�&���6������8�	��T��Vr7u���=�/��B�G���E�Ob��W�ͨC�#Ĝ���d�ɥZ-	�/�d����͗i��}���ͮ���lG�8��$eZS$�(^ �G۴��o��H8��$��h�{�̚����������#&Ǝa�X�� ϳsZ��ok�-�w�jD���o��q�>�QGךg�o�> ���f{�}�f�d"!��e{n���C�����IV e�w����ڛ�&M.M�_�d��/����<�y*�Ӱ��3b�n,��ո<0�a`i�ܶ�]Ρe �|����7Nk.��պ�&'^ޕ�5&є�O	��k���PxU��{�R��n�*�>�ÿm&�:�z���U�%�K�d�+�&�پo�)R��X�~;����]��GS��{���߄���Z�9lɆV@D�u��^���Ц���"��9��+�}O�����)��(p�����_��*p,�TTM*&���M��WuP���+:J/��ަ?��_t!Q�k@�v�&�O���r
߁[�G�(Y�AؤZ�|�].o�0&7�٘��^���W)��M�:آ5�����KII=Sg�|��fWTJLT��nW��P��j��R[@ʤ�hx#o�O��U�lٗ"GG2�3��!6bRL��Ŭה�?}�X�-H4�$%�R��ynמ�E%9�^BwZW|x��K=,=����;�zm(�ц��eXoX8�L���>��.��1�Ѕ����q���	�&DH����5`$��>I�$>�e]%OR���L%a�:�ѩZ%A�4��W#����]�8կI��v(f�8����������2�)Q�������qR�cF5�� �G53�@��נ$�3|J��ᱭ�}��]�n��x�_l��n�3H� �#�j�S�&�;N�V���nT����j_�g�Ļb��\�N<���Mj-�zWAf��(�ch���w�iP\,_L�.ٰ�9R�O̥gg�x����-<c����aaz~e(�"�6�������%:�LH���'eE���$ �Nx�	g"ؖ�����~�Հ�|��C�K���e��_s���`߷!ń��P�n3��p��G/�xc��kh���i?�+9��U��
j�7E;I,m�W�_���.��+J
��z����� Ϲ<홿�����|�����挗����5�=��_�����lzh;���낔���3��R���̠f-Y}�*s�ʂ��SJ�~��#j׎��|��>���u�=�t����i9��\�T�
�^\m;a�F�k�'�^��J����$�/tVZc����������\gߘF�v�I��v(�y9�6�A�/��ر�Q�����
QN��mRHXF��҂��H'�C�n�{�d2������nJ+g���'�q�&p����B���i��7�k*zs��66)|���{�BΈ��A�II��G�;��hsR�iС}$s:h�����&*)���o�y�1���u�OY��I=F���.�=�?[bn~&:�a
]���Bi;�`����'�t�`w�]n[V�ל�*��ԝNqQ��Doz���îaq���g����
�/�>�̝�a:�����أ#��{E�u��?ڍ�_����0�)��SE
<o-��⠋��;�=�F�����:8f, ..���c��!i��WY���̡[��.���g��;X0U�_���|~�̀I#y�.���p��"����4����+<^X��@ft�d|��
�UY�^=U��閭�3)��5��z:����#UY=����g�#��IH5��)�e�H���|@�>��!e|�o�F�	p.�����L�?���:HtƆ�C����[mR���C�@�-��¯�d���`���YK1i[�Ĵ�U9��9�4�.��s�H�P6�HV������δ���'g����V�$�(�R��|��-�X��!����p���at�rB��J����P�:�/Wa3=S����_~��R� �^�:W7���
��I��'g��9�9��K8�蓆��F�,���\��z�U�6(�H6����̿D�m�a����%�fh(���*����dbY_���xa������;u�0�鐉�M���nNk�9��g`!9OB��τĕ�9Vy\��\�.�d���ZW�3���6����[<P-m��/��;�f�D�6��&�	��$Eb�Փ���^��!�����8*�agm��anE��o�i���~��LEb�>ӱ���I�FA:��s�d
&�u�tT���1lW�����v��j/)j1֎�Y�
���L�<�:�(n���R��M��7`-�!��»��Uj�ቮ��d����Hc�f�����B��I���@�y����q��U�E��/�&��v�ɀ��H+D��i"!A��7b��$��c��b�����Y�eaw�ڠ3���9Q��S�(4�	� 6{��L��i�Ȣ5�Z(�����w�p����%W�{�lo�M���)�X����!}��:iaw�)���#�$z�p|$Z��B�\���Ԇ�ֵEk����m<��q� �b�{[o��:6���	���bIs�niiXڞ[�`�I�mL�����\܃�1U��n�0��D��������fd��{ �՚�)��Vv�OɛKu^>���I4���
�q���}��_-�e�?�a���o�e���n� J���Kb�����r�-�����>pD��ă�ύ$�!-�S����u��j��h��I���Z�i~��2E�Kìw��G�|�p6�-�6i�Y�2������B����(�����Ӟ�] ���Q�|xvj�pİ!!������� �WMA��F�x�E3���XM]��0	����dq��ؘ��{��w��{�;V����Wzќ-��T"���N��\#~�'\�C���VMeHڧгTC�]H������M����[�t.v��E��χw�>ɋ>]
SN�Rd�Ud�j��R�i���*��ϻasɊg�D�\��5W!��)X�?���l�s�[x��� �|MV_��h��i�!��>|k�C��­zyY6�|�MQ=^���J\�v���OzoYy�L��]��Xa�̂6>�0(r9�پ�	��7=���Ш�A��u���Ƶ)�Ԝ�ZuHHu0Ɲ�b����� �"��~9S&�s�R�U?U5$��gيD�w50��|.�2�:e������3�	�A/�-�b��'u2���i_��n��O�ת?� x-���w.N(څ���%JL9�v��Jh���#C3��eɎ5���Ůdu�ɫGf������M�:q��4A]>�n)�H�͠x(BN9�BOV���O�`sI�~��_}���)A
�ȉ�����g�J-��R�V+�EH�D6��S��J����v{O؎�Cp.B,fQ3�����'�`e�\<�n'ѵA���e��uY�a�{A	�I)�ƞ6fn	�Ӝ��G9�v��R#Z��E
)4�E��1s��b�R�6�%���u*s�TQ�+1��%��7�ד~_%��2�*b�v�/eAI�O����Y�۷�5bg�V�@���޳^ue�O�\�B�ݠ�;Z�en�js2P-^�dև�������U����g�;�V	��Ư�D��Z�7�no�^��"434�e�y��5��I|\G����()�)�%l!���\ASfb��v�#B�l���3�-�����h�#GV�PS� ��x#�d�3��<2� ����3�Сs��>��rÐ?-�U����j�
�,O�7*s���cQW9P��L�vrl?��mB��a���~P]p�>�r�N�#���������`4���n�ME��-T�&��x@3,ਉo<�|�HŌ?`[˸+9���\���Fރ��g���E�滟E����n�?�-7�R���߰5��D(Ń� �+�Z�#/e0��c$�~T�s�����Pm��߰*V�1k]y���;fiɽ��
&�8X�+���jC$�j����tg�����hB�L����F�`��G���+2��b��z���B<�RC�=E�pl��Nf����3�� 1�|���p��q�"޾��_E�|φ۔B����U����泻�v
ڶw]��2�=�I��D�ײ
�����Y�K��Y_�O�W��B�{�;H)����^n�<��DBh?)�Y��U�
Y7!ߖd�F�.��(s� 9i��*���g�h�A��N�^��RN	NYJ��'CC�����G
��n�nG�6�)���[1�R��������q#j��ȁZ%C�1�m
���x��e�I/� ��R��@�?s@��aG-�n88���%KtO�(���NS��D��)~�O&F��x�b�-ww�ceE 4Y�>m��ɵ�,xdcU�NQh�#1���^��ʢ����&r��(fq�9�gF�E�Z�82n�Ls3�����T�	Q�^�ś��L=ٽ��f����`[c��4��o)��c�=�Ĕ޶w�� އ���R h2h,�_�"!h��]�dcp	\�(�Y1���;/��7m@<z�i����	��D�����Y`�7��j���;��V�H斔��Ra����2�ԅm&�/	��/S�O��Hnv��#�PqF����3��v��2�`��4:�`�78W�&��u��K�e�n�s܇�r�o7���mdhQ���yo���xߦ�1b���,{�ɻQ��j@��ɜv�lI�A4��+�Xs,~����bR�f�5 ,���P<��Xh�6WVXV�
���g��OCл�m���z�%	���Ԩ�V��K��[Y�����5;���_�{V���#=f+?����~�;�H�ɾ	�����R�\;�&�R+�^�>kp���T��w���:��-`P