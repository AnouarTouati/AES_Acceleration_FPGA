��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&Ű��=�b��vT6�4��L�b,	/,A��"⽰k��b�t�u�zU ���� /��QU�:�4�S��\�r�q5�a�ۚN�PX�X��s,�I٨�iHĊ�w�����[R���Д6�N�1���_	�x~ѩŜ`��C���.ZV_W������K����#����Ԭw�% ��$rC�2��h��f�K+�"��kjҡ�V=	����v���%����*��*Z���o� *y�}B���:P����`T��L%S�n�����P9Q��,DMD $����4�P�� j�n-=�� �_�d3$���i�`�eIoG8;Z���<���
� v�a4�/5Qd��\56ù]�6�{~;��H�)x�П�q��y�j0��n�k3�2�S}�:���@K���`-��:h��#@^�p�����kW.+�� �X�~���������I���WgEsTg�z_�ؗD����M86)�c�U.���<�V�ݜ̐oek�1�/z��17�%�S��h9m/�By
a>�v�;e�_d=�����+�^塚�ߨ�B�3m���U�q�4�;
�r?�'5F-�Kr��Қ9��I'�G��nǦ�/�bT�Yzl���G]�[�_�^�tJ���s���<�#�ʀF`�JG����ny� �躰�_��t�J䧓Z�fh2�M{�F�?oxu;ô���>QmĢ��*')˪1�9�p����@B��&���'1�Ք���'�R5x�(it�%�� ��Z�-���^\�3���	_�x�����q{�-~��.�!�|��P[�$-� ���y3�� ����NMc��cW�iQ������\*���?N=I�1;�oρ��D�AYI�i�w�O~�gv�1���[\`9��<�G��M};������e �+T��Y�O�>�=El�����x�����=��C�[lJS��9n4Z?����`ħ��T=׾#3�cn�~�5P�D��KV�DH��ꓵ��7{�U�r+1UJ�˾H3��4�k(Ãle���u��5i�p�Xó%H������c�"�Ɏ��91ĔM
X��)�R�js]��C���5"�Ь�b<�"���gE����:w��Ԣ�֛��D�=� ������O-��\�f��W��v/��1���Þ�����&ͬ^ˑ�­�J��}h����l��)n�tD�7�r����9;�Y�����0�CD�sB̦�S)0[��.[�tE9���~�C�ӯ
9��Ǎ��Ӟ����^Z�p��Nh�V�NC�������i�ʵ��;~�6�e�>�v�:�zv|0y�G�Y9�4-B��#�X��̌�6^n���Jn��
H���< ���zq�����D�:|��E���e�lclu�#o�bç�ru��*D�`)���{�3�������D�(H���@��W��� �S��2�b�N��$H��o5�3�0���>`�)����e�����5~	E6Sb�Ҙ����k��NhS;z�B��g���vu˖��:�V	�$���U]��yI�֏xy�>�����r346v{{8N��IiG\�)n�g~��+�[)DIT7�ۮ�W*� ���i&�k��K����*|L=�+�5��}~�Ux����0C��m�,�O�a��#��`���Hϴ��z�-��{'�r�eh.O�4;�O��<�^.\>1���C�j�ǉUiQ��q�@h_������AG�Jj�5�d�Yl��$�D�Jog�S�C���gQ�V�1P�g�\��y)��گ��Ƞ�SK!rlk��2��{.��(�Ä��+f��n%�#���m}r���]%25�}	I������
β�rH��� ��;L�?Yn��$�^�������S�@�ں�Դ�P�Y�m԰Է=�ւ�˥�t�^��1gz�P�n,B޻�e����^;o���w�'�M+�D�4��񉸔ۿ�Jr���},!�1'�k��/���u��'��Nl`�k!ȥ\���m�Q���1u�]�r��Wp`>�����(�[�J��D�ѝ�E�!˚.{k�h���.�;�!��{蝺GP41J*bv�k�Y���+s�Ly$-���:��$e�H�Z�|8�bt
�|��;��gS5E�@���Q/�8)�|��I�ܑ>�@wɞp@�ŕ��@c�X�$��~ %u����"S��Y� �����',�"5B��2�t"�uÆWy)�R����{`�1�O�5��崔U�zJ�^�»�۶���B�~��Ib�b�D�}�x��B�F�0i�!<k�,%yj��N�Y��p�N��1�˥�Q����ۍ��-w�UĻ�^N1#6�je���~EejƦ�9+��3�*&�t��\�C=�y�_����mj�-�른~ �[0F�*F\�I-�ʟ�O������סS��v�'���kY'o�p��N���w�5-���$���r�ä_u�~MV|���iiH�#2�!˩��I& P�o�L��܏n������y+5����!�O~wH��b�+=�b�;׎Nj�ԁx��[���OΊ*����S�R��� l���Ӕ���`a��B.#�|bE�ϧ<	�1���:X�Xu��ք����WI�1k�����DׄxV4��Wt��J!� m`�-\d��tk���g#Y�Va�{m�}�}�b�ue��2���"��Q�Zk�8F�>���uc���w�������·}=�B�\�,v4��O����9������_��ܷ�;�0D��u:xI� �j>sG�|�d�!W*�
D���Q7���~5�#j�Qjw�4#�	���x�ygm6��;Z��;>8�~
�@�Ae��<G�ǩ�v�LɌ�-�O \�X������'�>bY�F��ZZ���ct���v?$��i��z��XF�c�}>�,�Un,Tj�S�(�<��0,��,0���� ��W+�/����t�/������ɻ����׮}l�5�%� �FIVf��{2�"�^��m�V�!l�ް\�SOC�TA��Є�%�5�bj�^��~��M�d	�|n��uW�"�qC�3�b,�P��Fm_g@���|��OߨE%W�FK��M��̒��vC�z�#'�&:6�7H�+��)��Gp8jsLT�%��8�Q�!> �J��G�D�v�r��1��0��c)S�"%�cܟ^(=�x�-�Ѵa��/m`�pk�M�a㬠 ;rv����6�����ۃ�p^C�3�6�=�*�u�=�)���۰H�i��/��N/Z�& Lۺ��z�K�vM�{Ou���l�`�'tn�~��`[˿��u(H-a��p��{� ZG�">��m|rV�� ����j,bb���q+eh�1�hUL��ϡ�G:�,�9��U,���M���j�G�,��6|T�w? t`�,�����uu��	[L�Zr��H-�O������_�W�b���,GbW5�S7ޜ�ҟ!��P��"�V80��]�]�⁒�MF�֥��4���8���uCQ�Td#��i� �����FK���/�����K;�zk�Ӆ�:fR�iG�kɑ��!@��Ew�:����Fyj���i��0�pr㦪u���m����af�/w��*\��.Z�T��5L��%-����?��NQ�M�TOuR�V0�%��^�dai�^i�v��`R�]KV��ŉ�]N�;��J���K�_��1k8V�2W��h@��L-Q���N���?s�H�)�%9�}(�q~4�sFJ�H�/K�|���=h\���'��kGx��/2�z�o�G|1���F�XM�&ڑAB9ݱ�
�}v�HG���-R�l� ��N���3�Gh6�x`�D��d%COy��3��ͧuy@�N?�[�.��c�t&:���͂��k[;���!m�bO�~�Y���A�T��s�V��%Y
Ÿ�F���N��kG���i�"R۷ �l��m�w�r%HcSM�O�^��F�%haܿ��Z�����B�
V!}=���e����w[�N�t�̛sde�V��y.������}Ooar����#�׽���? �<�/H�I�T�|Ǚ���}s�ҥ� Z�e�P��1�s��Om;r-�LY/���v�bF���>V*��~����VP<�йƜ���������� )bg[���;��[{6l��AҗG����į%'��i�a^�Ƨ�|�>%]��L4��rO�b|��Y��N�:�j/�����R��/���b�6��U��y9�s~2v��ۜ��/M��\�R����t�$/c��q��_���^��0��+NS��_O�ȴ|*�S~�3憽?	u�*b�pF�4�B�~IsH��bQD�>��.%c.�E��h2Wb�HQ=Y'?���۟��:YXs4@���K�d�a[L����y�(�Tg�`+Zt���i�v��bbh4�)�]mr����q�T�3+5�[��юH�%u*�IM5�F$ۀ�Bws��,�Ƹ��[{�G��h��W�$E�tJ��.`@Q>:V�_�eL�}�D���>��8�q��P���y|Ri���&��"s��z~���ѻ�qv�!���Ӳ>�R/C�&N|���M��D"��*�8B!� �шAg�ً��R@/]��&U� x^Ir��tǹ#�~����Ug������:4�P�\s;+.��]#�C�&� N��sQ=�T�z����_ ��1��e�$P�-?�!0�i�.Y�d�T4����.��p�|��C>�
}YH�C�Y���1�N"9���Q9��z���P}�v2�w4ҙ#v?���d�7�C9Qg:������mH�m2k��S\5�rK��������޸��۩
ub�xn��W�������f}��󻰈���\8���I�ʪM8�2m^ɜ���k��cW�@�p�]�L�q1�7ꗛ^�B��n�РUTc
m%�����\�Wz��"�-����@`�K9^%Az� +v�$�Ѥ�:�_���[`30q�ߧKdO�w�$�V��<3��.�#���:�nG>���u���R�0waR+ʄZf�,R��A~y��њ��0���`[WF���H�Tr*��K�I�/��,��
)�� ���1S�)N�J�$�:�?ZN3C `ka�fŧ[�\���0��ɣ}Y�[���p|Fq��2�����9���u���H��p'y4��������������l����n�׻��|/ �l"���(@�4�.�w�c�;<�)�?r2��u_OB
0�,���h(���n���	^�^��݈�{9�F`,J;N�z�d�?� �+��F�S3���I�4��L�tL=ִK+:�P��g�A��1ck41^����~����֛��5��.�RW����[`�qƓT�����:kM���l!�Oy�9��M�U��L�zH��(C-}��{<�{Z��s-��0�$b�[^��$�(Kk�zQ?���8R��xK&��Е�J�d��-ߢ2�	��nү��S���6K#�>Wi$�r�s@�A�h��(�]��pc�{��w��ot�5\=w@�&H��
*鵈AV�1�QY�l��<jє0UNH�tX��#�m���N�la͜��������E���Jh�DZ��,K���py�qZ3*h{/|��0G���S�癈ݘ"�i����x��w����=�j|��gU%w�Ǐ8�He	��4����~J��<9䵡��"ڜ�{���~Bl$5!6�f���G���Ȁ\��az_�ԇ�?Ƕ�*�7t�!�r�bZ����,���"����P�0���lE=��%n9��6*�NYq-׶ZLw���p �0�PgS�~#>�-�tWuF��W�a�7C����+�x��e#ٶ��уXN.���Բ2�d�4�N�g���b���%�C�M��)�e��ώM�0}�7+Rg�3J\s1LDi��zX�zA`�xD��6�n��C~0���8��	�^`�kϙ y<lɍ�d����F%�^c�"�X2�t�N?�U6�t#���~4WQ�'-5Q_�:��:p� $���_SOy[5KacYؕ��I��C�Lƈ]p����M�q�|�� 2���,7}��� ��;	��+ͫf[��w���#i{��o�=['����$N��܂[�� �K�^{"��+����J���v�
��1pr�����i�o0gk�ҙg0��ghN�jJK��N�𜿎�3�m)6ƈ�a.]۩!
�%ˈW��a��m���S}`MR�%g��A���<)�t�:�(����X�����{�^.���
�yP��������<�l�f��JM�Tܼ{�k�K���_;D/��ف�WJ�����o��SJ�Y��~���m�X:�L�"�v.��?�q��O�B��m��vP�B��p��8'��r���G|u3�>R{�S�uHo*��$H�Sy}YD�3��i8����^����#��Pa��e޿�f>�N��8�9"��͇l� ٥�"t�CM|����wfK8X��"��Q��#g.D@r��.�b�)hwF��S�T���^x�,�.@=�ؤ{<���ܪ@������mzgk�A||&��c9�=�$����=���vq��Y�D8�-@˺�\�%e��3�"���[��є�k�]�#�2��8�v?s�C�6?�	�:��������u0��}��R�5C
rF�}����{d�%�ϦUqI����@���έX	[���B��n+��=o����,��)Q,}��� ��x ��>�C�(8-�Vs}f�lUN#3���a���@�hߖ-�1��XG4
�D#:�.	��\X��T���B#�z�E�;�xH��[�[��҉�zs$=A�7D���-eA��i�tb~O�Eo�d��v=_཮#�H������f�)W�er���Ep)�4|�]]��5��}�Uk����/̖��іOb����fn�t:*.�c~��%HV������0RdZ�m�_���[��?��;q����v�T�Z���r<m�+�h ��ɣ�3C�WE�ݣ�b�Yv��G����_� 4���.�&�q~��,��MB#�D��o����I@l�.>�^�<��؅Нq�/�ѽU*�|am���4��y��[~ކ0�̎:A�_=��?O�+8���L�s���/h~T���ssX�aN����b�ؤ"�F���ڦ��5���U�LS�Cq�Қ? ],�D�8&�s`�J�U�fX��#��a�m����lcݫ�|�����5ol�m+�]	y�}
��c�	AG��N�A�Ni���"|�`^�ΔL�#�\M�'2�*�c�.����1������0�l����e9cۯ3|9�WE�A�_'�Mo�IPݧxpʼT���Fk��i����&:�Xɛ�� ��5�v@,&���E�e�����lȁ���ո�]�v�4������i��op�?^��~���(ba���
\0�I+�7|}�]�-:��g�;M]8�a:�Z.PG8��Ƌqn U���O�,$�^�&�%�!�f|թA��T�@{�1���(;�iR�u��2^�V�U
���
N+;�y3ӠZ�K�9�C��9�m�c�#�A�n���vi��ᝯ
��%4���T��e�)�ۗ�����7o�ϢI6�8��0$�w��<�
\�L��2+Ն?o�$f�l����A�����+��ӑzm�:,��Fco��=G�s�D="�L,U��S���"�q�hH����2K��.��)=B�E������̙^7�;�$�	ȉ�.�N�'{����5H�w�:�%l54�CR:qE����1�ڶ�׊��B���-�1~o@���}"�D��F@�����g9�h������5q�\V:�h� o�ub��&��=�2�-?�N�؏�a����Lc�lՏ�?^ی&��R����M|�.�Pfk �N��*'7��m�N��h ���y�LW<�ko�*.��8�P�O�Y�;��Q+����C�yK�!�?����g=B�t���:��<o�b�Q�^|)o��з-g�nc��}����iLEm�(l�5҂L���d�<�gX���I�amixG��bD�(�USx�� ��M�J	8Ů�G^��Qv����������+M؜�v�?����CLI���z�6�;��)��w�W��-Q�(�L|�����3n��'J$���7>�MSuU5)��^���H[��dx���/��ml��j�mL,�z�-���oә��9��{W_3_i�w�����+�<ws�>�#�-ZK�gl��+�g���Z�I�gC�l'��4��7k�"�� AT�1V���z��İ�0պ��̰�&NE�aȐ�� �*C�B_����P�$��^BԊYo
~�ֽ�z�������`�������R|a�mֳ;�;钛��}�K�Af2{��4i�/nӏ��/�p'���W��(\t �� ���
��W]Cu^E�56!5�E:굀e%�$���t�e�-�K���Y�-�j$h(l���!c������*�n@ Q���C�
�[�k��<�^U̼#iq�vB,��i��,ieY)4�3=+�5��]p��&�I�E����gP?�YS���/t�x+M�{�z�Z�\O6��~ȑJ��,}����@2�{���]�kYc��<�}�z�?��W�^)|�YF��S�G��A�Vrӆ(�>�qv��B�z�JlG�<����\�a�<e����DVR(����rԺ;%㋶�fF��R����ڲ������}��68���h�Z��C_��W��6�)� ��d#u'K)٥��r�o��+3�x�2Q��}0���;��x��DW0�Nܢ,�,� �,wX�m�	�δc%L�\�����P���f�x.�ެ;�3����
P>�?_��l����{�ӳңxOl�R��	X*�;af�A�s���g��+Mc��/�Y�(��3I:b\W��v�"Ę�~E�Nh�G	h��437bk���3�pͲ����^G?>'a��?q�ݣ�'�%B�Z�;��;#�!N��'�M�0�R�`��r�_a�5�7rt�%��,��Xp/j&t*(mzd}��,�j�!�B�F#%�l��U�=4�����_��]+�f�M��ou(�4�$�Vy���1��.:Ƕ��L}̞u}�s�V�̲e���k���Y�/�tN���vN��! #[/�K/��cU�)�v+���S���|����5�V���D�N�1_�<P+�b� ��?LJ7W���w8#A�äP���~������>XR�A����0���0��I�w^+sQ�֏�JXLU�@P�M�Ks�a�,�{��	�7�4�ޯ�s���w�!��BȔ*-1S)O��v�GIh)��J��7�����:~W�ݕ���c�Z��m�T��6,o-���������(h�l�J��L�뒨����f>�e���;�����8�W�a�t���٢��G���o%����،�ޡ�qo�_�"%:8 z����Ady�5�2��i˅n�b�\�Ƙ"��x�K<��+�ެ�)��r�pV=�oK`�H�%�����&�L�}��+�#����8�z���R�0�Y���u��*�@�q��slG����)b����^3���y,��E߲����f;��L?|bR@��˥P��n�K�,N��+F9����t]�ɻ:�aՑ���*�d�tg:6���+�ahM���M�����]��tZ���p �т�U��1y��ӖF@
[G���SDU^������N�Cj�<kĉ(��C�u�,�#�J����<����$^1�C�Xp��buS�1���|�=�\�D&��a>|q艍�8��;q�u/��s�F�8\�ϯʃ�Q�a�k�b������s�9;�+tO���okzi���' �at�Z��u&�߬�c��D�%L�ѵ�'��Y Ա֨*�,
����Ʊr-ٝ=��'�F�Z�$�iu�_ڎs�?}�K�4u��i<R�I�u_�V��u�x|�:{��ûs�G��W��!��`4�#N�4���N&It�[b4���-t=h�$:]�lu�3ǁ���Y-[�Ґ�r��\�^{��h\N�D�0�)3���ʃ��r��;�ߢ�}�� �@U;���{�M���T~Ǌ���:�PR��@�٢]o5�ęi#��^�u�ʘ�`py#�!�9���d�a^�9�*�6J=4N���p�@uq!�C�������f
k����Dk�!��ܐ�G@J�������-m��v��v��f@3ԛ�K!�9vd��A����`U�j�����>��>T�a��� u����f�� +�Gy���"�tS 4�j#M��	�P~">V�M�o�aX*o�
[��I�*2�b;���?����'|Bt@��N��g�dq�ԇ���,��hϱU����,�68���8��.(D�W� �'���}&�^[.��y~��� r�eKC���MF���3�/e�K#<|j�%i��"7�K�'l����������
��v����<��E���t�f���ScB�\L�}�7�6,�B6p��C��V���c�m��	>b�ť78�ڙClt*C�yv?@� O�]>@��?o��<��9yr-ʲw�b���c
���y]Q �0|%1�m���>7��2�4��z� ��
��,�E-��9�䃍���,0H7Z%���T�lb^+'Ρ�`�1�ue�~7��o��DL�����Hy)�h�d[>��%�{���v� ��o����ܓ�g��N Pw��?i���-._�ʁ��RQ��(�STW��]p��;r{3d5LѝeW��e���	a�U�JZ5pyC�:����MX��s�wx�Q����ٳa!l�*ʸ����d�/K�W>�x�'^�ʇ�͘���i�qJ�JI�2�5�4��1��ɫ�QJHo��[� $?A���˄��TE���ؘs�|�w$p�(u�Y��Q�h�&�E�܇�pl�r���tgE���"�jJJ,Ovh��1��d�g={�����w\��- �� �����>Rx�Եh�U\ձ�a��c�E��.����i 6����x'��+S����x�|������`ޓi�5� UV2T�z�_��K`3e:��������$��G	>#�'g�m�0�0���3�Y m�2�iQ>�����a6�=!iL6�C���C�T����m����xl����S�����k��M�Qq�Hk���W�{9�$V_��Ko��-���W���|[���������CAN���c�E ���/R�7�g���Vęs�%P����ك����$��I�g�iA/����2B�@�$�O�
�����;�T���$kծ{m�B#��$��_��{v���|��3Rz�w!�XF�����A�Z�HF�a�qY���I�"����C�M{mѿ�=�sh)�8�T���5<�"��TZ�p�V���h���,���RPj��{L=�j�6q�¤-�.��f�UL��o�"!S9Q�V�}����M#0�_�骀+|��Ҝ ;UV�S8K^�$��<s�z��+�,.=�Tq�W�r{��� F�W=�.b�W�4�ɞ�i`3�ɽ��\�*t��p��,�|����iW�܎˂"F���WWǇ0�]1B=�!�\�D��5a�RK�M���;+R5�4���N�-��r�#z�iq�I�;J��b6���ׅ`��eZ1m{ -#���/�+-T���7��`����:�����>�!K���3;yv�4a@d�;�X�_��k�T��P�d��-9'{�#�+F{D&f�b�h�d�5��f*_ֈ.�fy��`�Y�L��"���%���a3%����mL�#R��ErK����Q�t��Eh�oX�� N�z#^�z<��~l}�+���9��>�5���)��!���ծ��@d?�n�մ���� �9��t?=������cP@�(T)�������:eu�b�f���p̡�C���.��^+�Z�a>� I���!+���,g��m���˖{��ku����ى���k��j��OJ"�.b�l/�Էwc�]F]��m}�^�G�#W2J�o�T7f�½������)�݇������r.�RTm� ޵��˟L�� ��?��4�<��,�,�ľ��=N+.X�����c������(��B`��ۡz�,�߶�����G���(bIc���:�	�U�db�0L�C9�v~�޵U�}۠��L*4V[�w�I���.H�y\g1�t�:�F>(�!��l
������S�����]֒-[K�R�Pb�^6֨���0����W�(
<r?8�oT/��|'U7��)b���
�n`t���t�7�{n�.���w�+�ģ�3��5�W�zm"��^��Ǳ� /�r��)<^���q��O ���An�5�D�ĩ�KzƼ:N�#����cJ�'8?������b��f?�Ѭ�* �-�����a�߯6��vC^}Ҋ�|j-<��/ȺwY�6G��*�E[\���4��qv�t^8%���������[�G�R]�������@��|M��:̏/��}��eG�q�����b[��7"��m�Ob2���D�w���\-�M�lf�,����Sq���wgu,�F&�H1�>ƌk�@�rht���-�-�A��I��0Nx��9h�Rw6ٮ#K^4UECd�N��b7{-�%nI�x�Z�d�
�+"��K[9�](�>"us��5�(��g.e.��l�(�ϼ>]�$�ā]9H`З	C��E� �T�큳 �t�|��'TڢŜa��|��R�-#��I�9;lw=�_��O)g+��-���{����E2
Z �0.u����8��;IQ8Iؾ�C�MbZ�fW-˦�<U�?G�+~��✴�w)0'<����F���J�d'��JtÓ�Y}���D�[�z��g7yuM�D��h�ձ1�_�T�Q���8�D7�ln��\��2p4PH�����F���D8 8BG�T���p�d�|w�+bR8�!�����d�c�8� $KB*
��_x�n� �Yj�C5~ >GE��|e؀e��,���9LD�NQރ�=�A�Z���X�'��1�	����5�#��Mev�Ji�tE�G �P�~��\���aսh�oZ�h�o��׉�)���`�ς�a;�s��C<{�e]i�T����S�Y�-6GQ0���k{D�f�N[��YDe��&!��7a�n���-ƭ�Ϲm�@	��2��H8�T��<�R{d����7�5ʱ�͠�t��^Vc
����a�g:��B�P7�X9������H�v/m
ǷM>[6cMԙfx@4�^!���Y�aeRq��5���OY�1������/���s�vGR�ξ��H'fs�;�ۓ�L��i+QURakn��,���\e���h\�����|�rs�\4�����A��c��&���٬=���%~��pI��+�QOS��E4���^e;W��,k��#��ӕ猡��k\���/r��|�ٙ��)���PN.�Ff����8kY�;K����>��I��BG�1�Jဋ��X�,������XG�CoX8�*������DRy����~E �l9t(l���.l��o��R��Uf�V*�]G�%���In���-����v��a?��6+��[�޴�K�F�LH�� ���oZe}�5��'oTn���X8���;�v96������ЈE��]���L��dK7�g�.7=Xp�ϋc���.=�@=�F�շ~�y��D�g�;/��t�y�l�Īo=Yh������ӪTh�U��A~Z�~�A�S�Jԝ$Y4�wC��^�7"�\�/���P�/�w�z%�ko�>�X�9R|�.�dI1ڒdp��*W��`g����5��HI3�Ӝj{�m�l�a���C�&��f;���#$�x�6��p~N�C<��e����X��q����6��C2�������^�c����u�i])�vvG�j�z�Ƚ)����j�>�K�ɂ�pN��X=�e����v�E K=-�4�/�QvDE��j���6Jc=""�E�A������{�e�y�j�Y�.�u��? )���M��ݖ�>���H��dBό��o���c�s���u��-Fk ��Sr��O�Acd<���J�&_�է>Q����)�v�����G�Ŭ����O���(���$h��l����qw�F=�[���l�"�5Y�?���ۜ�C� 47��{��Yw�\��ŵ�KpO��݈�dG��M\��jWo�Ly�Q��Es4:�d���U�c�^����o�@|�£%������|�(*2��cʳ� ?Y�p�Pe�q��4�1�BC/Ҡl�۫g���Ƥ�Uu���B���J�����s,�;��Cs]^��p���#�;q�Q�J�t�u�ձ�ݩ~\�M���#�?'��I�{Sx���5��g���O�����GS+�.y4A��{>>e�<KV�s��}a��HIy�o���J�3iH��svex�J�i�8} ��$��$�&��݂%�Bjm�/����Lru4�9>�?������$���$����'ЏAq����pn){cY�E�{j8�no�*��VjR=N�Y�\�w���Q(�%�DQ[+D�.�7�DW}�����nҝ	OA�C�T�0�-_G��C��]Ti�8����� ����]y��_�P0�p�����5�3+�@
���}3l���?t���U�ɠ��k�0otc+���X8͛u�]�T�t��Vf��=�*���c�M���z���� 2��#�"1o�|M���i�B
�����h*]�*��q�('O�h�3��+���|M���̸��7+>��KǠjkJ��pq+���.�cm�.~.	c��Zպ~GA�h'CB�G�_$�a�8�!U�b��T��6l�4:�˛������BSڈ�����D+oŀ����	�jF�j��W{E4>hӦm�����(Uݐ���`��a��c/����%Ų;�BDo���yiO�+�K�]y���5���?;�W���p,*��9oS+�y.3�mf�s",�z�Oc_�g�9_@���g&P�~�u��%.Z|�#��P���
��]5+�lt�R�AO&��lo%g���ܺ����oQ�a��z�O�����c��lF��yu�'��7�e?_�S��Y���,'�u��*@>�tl���ԛ�U��k��'�<�7��߽ZYq�v��1�9� ++x ��&!u���r_��,���@�,��䥉��U!��i�q��ymRQT��EFg���b��ܸT䭈�1�K����/�nuq��0W�Ci:�,h5H�;\Z��jZs ڪ 0w�i;�g`��.7l|�c<�#D6E��"�T�97E�]��5�Zx{\��ϻ�ʏ[5�vFugqf:U��q	9�4�6���ivG�gm��@qc�3]���y~wI��8��Z���.��P��^����+��H���|��Hݯ.�\�9���e���3-ކ�տ�A����}���2���[Φ	�����$U����i��V3?�C��9�Ȟ�Y� ��;X�Z�I��#R�,� ��7BG�W�ޙV|���v�]�ֳe��#ߊE��W���ɞ,���Jd���sb�.�H;{�54]��9T}V��(�`�h慓Fg�w�a�g&Ŗ��xs� �U�ext6$��; =�������,�:i�5�d�H0�褰�V,47���B~i9V�'�'�a�Q���>�C1ǯ(A��\r:#�^����q����FF`e^㗃 ~�g��_/��~N-֔����9�䉚_���
넳����{��O���'�l��g' ��w�� �2n�x�����6S��I.$s=0�*CW.#3��?�\5� T�@|smj��d�攡��Uَ?L��j՞$�ʲ_t�/-{��R�z��+�������s[b��.]�?ۡ<
S�u%vƉ��,+��($UzEb�L$�@��7��u=��Ì�Wd�R�u{�c!K�Z�)�T��`�!�� S�#�)e��W����,�s�TK�E���[��Vp�+�о���{�i����f�Z49��+e�7��p�i���3䞰�7���H)9oY~O�4��]�l�8������sV����	���KޱL��hR)�p�J�t�,�d��^���p��M5��Om9��t�[��MNю���=z��޽��2_��/%�"մ�P���u16�Fom�h��D������t4%����L�� �Al��w��_#M���'�38,����bD�%5�B��"I��u�89T����0�ҟ%���J<�H<���]���h�}�t�O&^s�IQŮ���t��RZ���_�r~�G{�\���'��n3��@K�|(�l��I�C�K/�9�9ǋ��{��Т�(��ǔw��@ԉ�H�����h$���k�NG���2����uÂK �S(�M���v�|�"N�Hp�0e1���;$��J�e�����i���h�Ƿ��k�/6��Ԛ��M7;�D�k&l��l����2Nrݦe�d �B品���(]�rW��-X���|�m9�,�K�8�Q��Nr׀��z��ǣ�$�����h��<q#��f/��XcKw��Yd��u��>'S�y�~9M`�5���:iH��ӕ���f�NtM�Ȓ���R��.;ǜ�3�/O!Vn��Q.a ���V �vtg���!nS­;AU��҅jSz�.��lB�G�$�`+#��#2����8����8:|B�|�ަD�O�4�����f�	nl���3o��2�d5�vf��W3T�:�L"�	��ȗ�=����Γk�l��duQ7��'m������J5�F\�������3�ͥ�oxS�YD�
�i�� ���^Ĳy��]v�4E���vF7�g�A�:\�U�
��s���0ѐ������M�A�1��+��߂���$�-r�U��!�̤Uo:_{ o�<պ��]���U�ϓ�"���*���zrWuT�ʚ8Gg{�F�sE�	G2�k(�T.�x)�(d�ܝ�������´�Q�Q�{ ���T�Ehv�\�w$�U��O�o�<Г)�l��8G��;�� {�����j��V�̬�?ӗõ4,:�8{��u�|H�w*��$�18��F��B��^�}Rf.T�%�k�?��6������pW�IN���zA/~:�tu���#�Y˒�B$��ue�jf����&m���{���/h�Sـ�����7�}\v5#��'���u5���':U��%-T��P�f3$��R�k�gV����nČ�x�ugHդ���d
bx�H���/��0��(T��*R�l7�������m�vu���S?�.��.�~1Yzg����GŢ0:�b%|�[���L�U\�7tP6D����� �,O��U�����Wv��%�^�準�>N�b��<���s�'F�jI�}�Rx�;��ʣ�,QĠ-X5�����7�Z/�>ㅳ���.Z��Sbk�~��y�
�M?��f���C�
�(��5���a;?�SQx\Qh�;��X*�ԟ��^&�t,p(��A�~�?�b� 9}<o���V_�\~C��9�'Hɥb>|_�\ħj��8$
F�t 0QW�����Tj.�6��(��i��}�'T�l�����ݸ���3EǤ�s)��W�F;9:!�"�$,���|;��Dj��� �f��|u�+�������27'5����.����΂��V�(azs�l���1�V�7�3����)�?�sNR��#Y��a��4Y���m#�{ �)��B�T���7
M=����t�V{~%�Կ��*�.>��6���-�N*�۝F�����#;m ��ׯ�m"8��\ڿB�B#����G���M� ��an)��'�ۑ�~�`�Sڍi��S���/;�tX�O���}ؖѨ]:���Q���8?*�h�;2�6�v�윫���8=��Q���.1���hi�E������9���B~�BM�冨��������<�z����熽mI������� c���#$!��U>��ٸ�{k��R� �s�p�Ir^V���d×M����� Yf�
g8�.�x������A�Q��NF'w�zk���궭�����.�퍯���	�[�$�<QD7O��x�9<�ǎD������@-�.��O�V8��Ǯͻ�C&�.Q.��i���4%
%U�>#<�Mc� ���Rm���j�Lj���;��z�-�o\���i�3C�r�R��V���Y��*������9�T�gi�=����"����F�gy	�q�x�Nj)�w��I�a�457zW	��
�?����|��F}�����8����G���w��`:�x�56���"��xo߰[�xg��>Z?���$H�N+qk}�5�6���t��Ԙ��nB8�Q���x��Y@w��т0_��	�����h>�f Bп�"	�#�n�����\���hcf:`��oͣ�Y��G�����n֕
�oO_��w�<�4��t�9�]-I,eǏǘ~���;�$r@4���^��?P��jn���xX���˰X��˾x�n�E^ bXr($������~�����Z��x��'q��;�ā,�
��γOڑk���?��d�O�62,ح]a��C0=��{�FW�Э����yE�
�i�����ݣ�O�(S	"
[7_�~Y�u8��`M�������i���Xv��KC�L������@�.g����^�5o��jm���]Ub�&�>�-E,��A�# |�3}=ԡeM��<�)��o�#��E��mzG����|]��
��9�낯�!����&�9�9�m�]��D���ʊ��Lq�J=wA��`���
>K���t���n4�ymT��d�VU*�C�g���L��d�z��k�<�@��UǨ�)�;8Q,c�2��u4����H0�G���0�M��}D�#F�������g��X���0۰�"����FC;��dB�D��
_�?�ވcV�n���(�Uٰ ���۽��s�S,B󧣉0�pXw��Z�v;씶�7&�ZA��9�ͧQ��N��k�З��i��IM�L~]H�No��<b�̎���#��A���2��=pA�_�i�Pa����&AU�H�-+�6�*�U3f�^�GO�Nf[΄/����&�5��!*v���H������1�IJY��h7>w��^c���7�0f�J���o�'!nd���x����bd��NQ�$�y�`n�&r�����2��QaFE� �OnA/@���gV4�`j�Ce,����xl�;��*��G��H�(!	/��գc1!�Cbؐ��^Ձ���_T6%�7��i�xd����D���+�3族?�T5~�\��v� ߲a8��mS�V	�WL�[��=
�=�6�������IP�Z�9�����g} v!�7���i<a�+�ß��t�o�����s yCOO�ϯ��&�L)7�������~�=����Wkct@MI��m�.�]��H���U҄q�u��M�8���b"��|����|�c`%O���mM�w��.�-/�Iy��u�|��,�|�\>�j����"����M��B.���ڲ�0��G�����Pݽ]�F�п�1��3~)�0i����)]U��+to�yK�@oܫAhzK�E�)gn�Tq����j��a��4�����B0-�\Vƒ��'Z}���	���m��ߊ �q�[c� �A����Ʒ�o�v� YƖ�Zsi�F�ƶ����<T"��Q�,�ֈ%�n;7���x!p��B6��v��vl1�CCfl�b
YM���9͸�/Ȅ"߹Ij�C����R��������e܋?�`�˩;�����S�)�����0a�ٛ���A�ٯT������N�WڐI4m���k���\���E�1oe��'�Ah5���{��x��	���S���K@7c�X�B=�r-���wҀ*��fy���E>���:�bs���k�g�����r��r���'��zi�t�	���<;�=�"{�o
����=�.�	�|���;���GYv0|��i�
5>)��{�vQX;��c���G|�M����V�W�C�
�Z�I��E�B�z�j;��h��F��*�ҩz.��9���R�`��{�%Md���uKI���t �7;at�z⺼,kM[F�~Y(B����PE�	��3oG�9߇�s��$	pp�*K�l�W^��X�˘�&`D��tf��w�A��E��A�i!�0\���P�����8�:�%$����A�fRH���Q�y�
���8�o�F�b����5r��"���ծCF�
 ���Q��/ꅟÇc �q�+lX-��>��%9��D�y����� AedY�gȱ)�V�W'����j�TB���񥍎L��Z��ւ�#Ѹ:�̞~�3��q�0A����j�J�KƎ����a���5C��zBJ�:�\8�Á�+zf��$�Ơ��{�a��z ���qw���&��ؚS�_��+��ي![_��H|Y��f["A�q��8���Jb{Y��b	/�?���tTu���� �8�)�Ќ�:�5�gD`���'ćO�y��m����	����2�����ruպ�������Q��O?�YR���Dh�����w=�t�4ܘh:;, s�L�%���Ś@�_bL^����Q������G��j_y����6[���C�o���� 5�)�]O�gF��1[uՙ�f��cO|׬��z.���TU��T���C��%�.��b:�i>�8OrKhL��6II����D�nZW�y߉
�CB�qbx��\ڦ;0E�����D�p،a���I�/u�k)\��~�$�U�L:���O���d�RjF�O����T�mz���X�p�\��	PQ��vs�sﵜ�A��Q��x��ձ��$��_{��Gur�2]�������(1�x�6D
[����u:���LWA�4}�:���i%��,��	�^�cT{�Qq����˃�M"�/�A�G>J�cڈ�R<�M �Y�4}���)U�(IÇ�j��MG���`��T�rX���R�R�p�~�Λ�b��i�������/Pdu���K>�?Z������%g�H\,ȋ���`�STSD]�2�K�����1~��u��4�ϛ�(нy˩G�6�7^8��d����������gv��({�̗;�f��(���QY�	���ymY�5v�;*ԑ��0��k�?]�͏b���%���O^��1�k��
�zP,�..���*73�� �*'�L�� �b|���K�ͦc�X1�����_V8�w�y�g1��E������d�70H�I��I�7GI9���s.)�uVoE�؎�o��
$Y���`���5j�SD�;sR	÷��̉��Đ��4���0d_�=��x�a\� ���K���PUN:ZX�c��E�s\��q�IT"�2�3�c\��biZ��"?�7P��Ϩ������C�"��� � ��fz4��V?�L��������'htb&r����dG���Zߞ�BO����'���<U���<�.я���V� �QTuT�zۀ���gxs�D����b�c��;�`��{�a�R���:ϰt�͒'[b��`}��ף�68�9��O�KI�/�k�@��up�5ֈ�)����O��%�A��me���R;��ۧp��& �秐�-��a,8�P�e����n�ga���Д3�&���r�g����1�W~�_����S�M���ݼ9��iқW��g�L�6.՜��Yvm*za/Ձ��7#�~e�>��Xe�A�[�"�o�(�Q
�G6|��a�E�����xo٩�n�̚nIh7�
����]?ѻr����{-�;��쟹d���)���v� J�U���-j���!����Wh:��]2Q��e�D�߲�H!�g3���҉bǀ�B`*�;���6^O/=⨨�p�Ӹ7�i����_��s���mNck!9>y�:������+Z��ɳ���T��uݱ��e٦1�X���j��Xd�D��%�#/��\��)�>}ρ�T	�-A�cf%K�ڹb�?�ѕ)�L6P�����x�����Z
}����`sYd�+�wY	(nYЬ�&���sZ�̦b�P�x���t�4��d3W��l��^��O�(��~�ޛ�ڣ�|� @��8u���Q��.;�9�º�� �l�+�/�m�Q6�-�A0����BU��A�