��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�oA��J�O3�3�l�_��m����G��ml_��:�Xc��<BQ���w~+6 ����[c�Ox�	�Cd���G��S�,/lY ���8��F6T���-�j_�0���X�&�)o��Ѿ?J�)Bxr�T��i|&�
]w�V��.D�'��XX1��A_T<ڛ˹�P��IT�`���������+D�}�c%�����9��/�c<L"v�X�&���o|2.���%r���-`����&�~���޵G2�7J���l;�����H�b�~�@ �\�*�`c�ɭl�? �B�B,��b����i���7�5V����V����᠌��ޚ#�P�Ѱ�� p�[D
��n]e��K?� 
+*��Ė�jH���X��������-��(���Ja[���<~>�q6GsO���hf!�p���D��O�|���G��T�_��Ƣ�R��!޼����8nT+�J��\o(��l��釢)����Ց��ְ�s��_Vg��T9�@N����#+#Ê��M3��V�|���#�Lz"�Ws��ӝ�us)�s&Ƃ�B9}��)�����K?��M޺�Ӯ$��[Y��;�=��+��3�#�}�o=��3	@����z��^	� ���	����>��+�jɵ<E�?����N-Pu�4h�|'��U�f�R�v)��2F��.��,a�\EL�l���n7S���D{7�䟏��O�'���D2�X9{?Z%���ts��ҷҁ�ݜ����r�������w�i�/4�i�`C����J��i� ��
C�ݡ!�G�p����>`Am�7D�4�a�Z����ɳ�af���L�XҜ�GW�����ev��i���S}�������>�W=�����c&:�P�t�R�����&x���t� ,����^
a>�:2�N]57~mOJlH�/���?�<��Q���\p:	�sf��=_gw$�}�Z=�|H��2m9��K�x]h�E`M��\�R
�n9�Fϳ����Ĉe��j��ʁ@�a��p���5���&s�s���2OOH�iրw�q�VF����SkL�22L�����/�����q��#�V�5�f���ѶO!U�ah�"wj�V����1���ħ�/�ٳ��o��ך�y�.�,V>1IG�r�=ZT�J�P ��G��<��-e����Ӆ��KJi��� ���1s�a��K��Y�k���I81�ف�������]��9?	#��C��l�4w�͘kH�36C9��u�zv��k�Qdm�v�������M"m�j.ܕ���qw����G")��xh�qǬO���4q1I���`:�_z�3��Qۻ�
�X
jgEˋt���䷊�0n�2 )%6��~��Y��1����K1�)��l+�2h�����	a��$��Հ��Ҡr��M-?���8m��~(���5����^e?L�v�b1�i�/�]��_����rJ�����7L�ʜ?��o2�z�k�kI��=~`�
�ӋW2��8j�����C0�3���#������e�����:�U�U�,9��D�c:x�JfGRy�.�\�v����r���,p�Ð^-:3L
Z���3ײP������ʺ�9 w��[���COFt�l�M���V�X���Z�6Q��-�r�v T<�n��Q�'���k�Uz�i�Za���Z�"?�9��N��N��9#�Z�.��M�6*�Ia@R����;�g��ѹ�M���.��Z����ǢK=��jQ������^�b*���j'����E��P,v&��޶Z۬{A�ڋ��A1Q�m:#2�ԋ��g/���G ݧk~W&���+p1kR����f�,<��5K�����V^0�LBm��?�r�1|�F��m��T����]��i5w�T�:�
GR&<�iK-�3�I��|k�S.C�=�J�q+_z����-�:��ߌ
^�o�d9iOɉNj�,X���������Ճ�R��F�dk�D �8��lx����&�M�3j�w9�C˂<�J����=$.[;�&7C�QήM���}]h�$�mR�nd�g��0@�a�;��L<��=���VbT0kO���q�Q���/lfB�0ѭ�Sz�k�a�l����5JN�r�]�P����f\��/H�@K��W>�p�G�칳-�6:��.���y�a��2j�{6��w�:m7���FNU�B����"U55rD�Gޑ��k"ǃݑ��/b:���]dm1w�п`#�쮱��;s�d�_>��Til"*���z�|$P��.=�\�1�270W�q��l_c.3��]n��۷P2�dھ};�M�+>$7���, >N�3rB�ۑV�E�W��]Z����a�6�ǖ�J�[�3���ǰ'���y�^4��O��W���j?궛c����������y�P���c�Ak��b��B�r|����+�5�������+�ˉKK��%��f]���p2D���]���#��0�����A�:�Ni��S.�BpIH q3^�i�G&΀Ȟ����#/�0���@�T���\��A�G��
�fRu^����q�)P����7���σy49�+�$��d��mZ���N
~���,g��2��*wG@f R�ݫ�~p���Pi������j��	�SRp"�˸^ \x�?/�+����J�5��H���SDS+95��c�s��mz�Qi"%�7%g�2�8�����!2�#͙R_i���q2t����6z��K��?�(.zZ�&���b��	M�Y@�(�5�������aY�U��#	 /�
蒣e�{����x5����������]�����
�q�lF9�����I��p}K}���U�x&C������@��i� ?���ݞ�����E$u���RZ�=���3x9�*_�_.� US O�ё�J�@'��*�D)V��3��k�v �v��8�IHS6,��U����ǍI�M��꜇O��SS�
��b!EI)�#ҍ�+�`��¸YO����d���O� I��������[D����M /Ӿ�v�"E�l���7�3x �����6�|	�\�_��}��BOX✼�L���0:���(�7�GwU�%�U�x�Ay]��ۑ1$>=6ź�c8Vǚ��~{:���D���N�F�ʂ�TuL��6N��Iϩ,�{�		7��|��*�=Z��,�kq:I��ׄ��:<�j��k2�0�
 ~�N�b���#�R3��#����[h5�K	�/
b�T�a�P�RG���+)�U� �'P^��	����}��R��(�(���<����	�� ��t��q0s���>��ݩi���m4��(�%�F��(ݳs���^Ĕ�Nu�p���f]&]��>:�y&Ң]��]�,����q\q6s�Ts�*V�م�l�Ť�顂��s)o9�����P��M��v2�:�g���F��DD�&�H3G�x�>t�3A�ق�R;�^�1e���u(B���~�tB^VF����+�OFX�t0�Q�z��y#�7E�˽ާ���i:�m�G�S.Ն ˸!���â�6��j�ʘ�T��`����N�a$$�M��L�\#���[$5'��g��ш�^"��9�t6+�42��ͪ��׬B(-�w ���2ּ���K�� �%u^�J�O���A��.��p�^e�m5�u,��?�t��JS#.�%�e�}n���ّ<��x �m%��P��d������s|�f�]�,w�����Bu�dt�UʗI�N�l��<�\=�`{�a�`*��)��%��L��RD4\L�/�L����i'��VI���$�����(�������<l������[I)�=rm.�Q��%�F�<�WS�_@XZl\��gH�f���=^6ӟA}���3��PGc^�R��c9�h���r�f�#o�����2��r2*m/������H�EG�K{�x:��{�	�?f�S�
�څ���^nr��08)|�6������3���KR/h�LUrw��n�bcl[\x�V��q>d������"���#��6H�4.�i�S���ZK�3Nb4=;t&��[?1ɡƲ^}XR6�!*f����O;ق�䐑�T���+�c�����然�s�*U���/&s���e�+�{�����OoJ�nB��`������$����A3���?e��^��&	x���(B�~���o�NQ�� ��*[��41�1��.���ۄ �[$��=*�
�vv���a�0PU ��DN�^3���M��-�X�J����������S�����.�
(Kd,Z<B��"�K�;ZV���Q�yXw�y&3�J����NgS�Zt�؈̆4 i[M���F��,�^�������' '�c\6J���8L�'_����dc.W]}z�ag&�(='lu)�O�=.i�`=Qm�3�I��fJ���^�b�	����葘�X�UZE�*��e[t�48�F9��1�<����a3���(��	�}=V'x�5oQ����}�U����g�2:��:ƍ5�'ɤ%Y�'�0s�E�|���̹�@oҢ�`D�����o���w�bh� !Z��U�a2�fWŧl�c>��	_>oNݷү+�	9�LQ"�x�w�b��~� �Ȩ~�����!S���ˉ�Af.8�W���x��:A��9B���~�N̴�-�-��/m-l�����e'�H��(�?ڶh+�r��f�D�:�/�;;��۷��CxW`Q�4>Lk;V�g8���4d8��"��[W��J�n<	������ed�CG.���4��`�L��EJG�U�ZO�c�{�k��|/��aC�;�</�C�x�'��*`�9:\�_Z܌���WR���Ehx�L9[�4 �ӟB+��~���ͻ�p������-5������[��s2"R��oq�J�8�~��H��z����ҝ����9�G��Vׇ���NC^=��3>?8�[�9���,1��q�r~�)��m��]tap�z-�C:�
�S��wu�}#_#���e�E}C'N��Δa	[�w.k�@���I�Q{d�c��`��9G�Zr�|�F,2t�A����F�����@�U9ԃ��Ei��&�ߡ�VW��[��}SlA�x |%�:�nަ`�2zڷ�	�O��� �Q0��[�3Y�ps]��j�Sv3�?o�'��Gr��r<�TO�+uV�uwm/u�9<��`$����}\p�(nA�Eݬ�`�E32��h������_����kR� ^;�����#=I�tE��u���ԩ�������+2�|�#u�9����[��D�"]��5��6ηygs��ǵ��������y�F�T*5���I�ڽ'�ju�����L�M4�Bf_ł�ۭ0�gɋ+g����M�<�$�GT� ��ڨ>`^K1�J3�����8�g��(�3��(n��Q�Q�����, B�-e��BӜfY`��n��$.�c�c��2Ղ߲�ݳп,؉�_��b�"������rK���j�s��&�J�s,�� �+�H.�Buw�����w: ��V|֏���-���/��cS����9eHn2�*+�ӯ˱�5t(`a!Ի'-��VN���S��oz�5� �P<�Ȇ��V�}t��e��?�R�)�1O��Y��9���ؕhP�Vx�z�H��g��K ����&ջ�_,��,�R,�֎N���0.�@Ks��U4X2=x}�ҁ4�� �4u�}����������>�V��	*�d��T�?E��gP"��s�o�qN�o%��u#�$OqE�t��Vd�),;�c���⻸vJƖ�@� c�������w��j$?ѦgT.-��n`V��<�>���{۝�O�	��8h��	-@�-�2�����2�O�#�	�$Os �*�?pP���qʩ�I(.lG��i5���ryA�Z�V�ܵ�0fa�.��-��]����W�����&��lϼ�o��W��?`��C+�7��
�-� HO�#�r���[�s/�׮�f�N���W�/����+��e��E���Y�%/K��D���H��S3Yn����}J��["G���#M`��l��+�?<�;��B�$�;�B`��ĝ%̳�����'�ӵV��75����&�Y��16�v~�Wl|h��N�]��FL�>���#��aW�AI:m��kos�T�xX��`���%��a5(�G|�&26�&	&������L���$�'�!mi�Q�w�����Ӄ�\��]�����F҄}����t�*|5��������4�7��ݥys9?�(L@�@��B���P%��BH^Ɓ��ae��s�R�DTq��=D-vƟ����G�9�aY������-�p}6\Ɉ��ـ�:���[��E�H��e�"Ho��׬%�9�mܞ��C��#]��eÈ�Y���LN4��|OSx�E�{��R�Z⥱.6�d���0�ήx��r@������9!DR匓.V��h�{0�u>ǐ�H���}�=�]DW�_���5?�Br��I�Y�L�� qo��W��J1S��"4���N��g)]|0�%b���=�ǂ��W������V:f*�[+�^���`��B���թ_U�I���v* �c���_�r4�u_�^�SUw��@R�k����
j����-"�����W p!���`̧<�����ܑ+�6�mW{�1+�X��<%���KY:HV�f��9V1�+?u�SPj.Ѫ]| �w{�U����,�ʾ+��ߊSW�ީLx�kW�>b�,�ܑ�3�X��SS$��T�]�Z��$L�6�hF�8Rrqŧ�Cz�K�&�W���
(#�F�q�-����bB�9��/iRT���~:y� _`�a
9�%���y�5�8�ѥ��O�֯M���H
I�"of�E�-�K6!�r���g��P	՟`K5ꋯ˛��;+�t��}r��'^���r:��lMr,�&w���pb�@r,^��
�p|��8e���;���ܘ�Ul��i��W:s����$,�Z�J��K�i��8����C�
�K�	;����fz`��bkԆ��ٜ�C��X^l�M����o�  ����.�z�)$	p�o�Fc�����2�~�������I{F�]ڟ{���ɉu<��Kۃ�z�M� R@�R����2�e�7�޸����"(���4�
��o���4;�_ �A+�i���Np:���E�����9�qOq"�tp���Q�vO��\+md����p�/,���#/U�p�d��LQ��!�os�dH�覺��3�ME׭ �����%��T�u�QEo�X�ɗ��Q���02Gb|���%�{����+w���-� ���FD��W�-��>�钧�EE,���^�ǌ�sq��R��a�$���N��b�L�&D^�CU��bH[/~��#���mh��`?��l��8�"0j&p��w�ݺ�SmA�..sV��|(H������٧��ǥ���}*iN}ˤ<���ޱ3ի��w*��#5���l�|��ΐ>���a�=Q���40l!%��,�R3��<QK-��ֺ 3+�K��@���Q��\�t�����5['ZwsG��R�)0�ݣm+"Z�'�ҵ-p~����G�=���=Ds�˙��Z�-�`�S��]��꾥�bMf�%*!��T��7�M��Jw���D���}���'�$�~6g4�/A_�K�h�ˆp�Yfr�ۯ��v�~�<����b�{
�0[k�I���Q_���s�=KnC�p��I~S�~�������D��y��������J�3[�X��5��:�x�1���f��2	 �w�({kt%J>�e�e|��
Lpk��/�c7�.f�E_= ����Q��B˙L.�����Z��wK.��5�J�B�4n�Z�	Q3��ZӪDM��s�l���A�Q�8�VK�8� ��wή��ݷ�t~*~`��?W�� �Φ�\\����:��۝��pj�B9j�Ff��ؚ�&(P����'3� $χ5n�Rj�������|{+ķ7��&<��db���X��|�)ƅzI62@��� ����>��owz*A�fc�y���#É��x��80s}t(�J�0�S��cB�E�j+P��,�� Ր|�6D�ڽ]4r�.��T/b�mrv:n�;OB����� ������y��v�K2�2ws�	���KˬqC����ƽ�
�hM�^�=�gd�3#=g&��U��������2��R�ze�Sx����:�FE%�_ג�$X̴ �۫ UxGbh��j#q���/A��[yC�&᜕y��ʷػ�)]s��#o�r���b`ouQ���^>=>��;Nd*k���h�WoFkh4�i ��D��d!��N���+_EG?Ĝ�N�oE��Q��}u��<�O{�_�3à�wy5�~��!1�j�K�
~UIjd��J��F�N�!����#?I����3��s�O�.�n�������sxC�UNO���\�=
��t���d�N��nU�-?t��S�����0΋������ҨA�Z���-F�k�;AE���u��)�����a�A�(��R���V�3���4���=��)K��z��,��3K�{��k��/4�x%�����zd���f1jX���?"��1+5�х.���Ep�o�pӻQKy�q�c�����6�!��N9C�����~�>@6�)��ߓ���Ax�-��z��1�X�;�υC�;�����ٮ�s:�VVn�� e�?�a#ZRa�-��QW �\�\4u��)���+��f��$����ؾ�xf���e{�(^��S TŜ!r��6Q�]�[�)��J���&N�j����e�ƶ���{eY���Ol֎,G���J���(�v��j�Z���=͏�
Ts��W#C�FO���V�@M�lZk�?���_�^W������+��F~7|��䃒��)���%/:�� �$��v��Ȏ|�,x��_ ܌��QkG�?��ݑ[<;qI$����t �F!���6�\b����hM�p��$�oः�a[��j���oD�Y�k!r��U��F���8ס�/� �(�r��6��:r�4�).��;aM��aN������D����[��2Y�̮�?��uYO�67��7�QN���se��Ǔ5a]�e�8<t��U����FxW�	/��d�QR���k��걑�n�L��[�,����M�c�O�����a�s@W��Mf; ߅1h#�iɞd�����yuhcČ�`Ad\_�������l!���JR�O�e��B�6[�uGٳ�P� %�Lh�?~��yK2���)�7�nU��%O�b��=�`<�Ũҗ�=�R8oBr�ٷM��~ �Ρ]�U����^�?�;ȉ3ؒ�P_`�(~��M�)oG�2�Yt�2	~h�g�~�7�<.���,[��]	�D�g(��ü�L:/̼�ҡ��0�]y�\L���/p��l��~���0`ׅip5}ӫ��S+4>buf�v����N;�*�bw��q�feޣ1D6]]�|x#�ֱ��)ߤ�H�z��^D�BԸe����2/�Z�Fx����U�Ω������g��[�T�d�`��ҷ��Sv'�]Nf�CP|3��u�a��(��~�Bww7Ż�����܌��G�hl�� �̳�'A]���}��I�⾱�t�H��t��z%�W�&�Xu��B��BR����^���j����8�C`�pk%(��X�⟿~�9����~��D����
+T@���H��p/�U+�ȝ�a���PM:"'�ᡱ�|q
Z&�Pc�v"�ǎU����/Wb�#B�U�pUɽjM�t=�DZ����yG�,٦QZ�fŌ/���*4���XH=�;��g�WF��z��]f�)5��Euh�M6c���kE�I>��_����|q ��\�D8j>�,$���	��u,�}�+7��գ���7���sx�[��헪���޶z���}��C]'.��lo�����OX��z+��n�V#���FD�R��
E�OK��n6��ڜE sz��}�p�1�s�fMW�xz9�E 扟Ee�h�2)��}��x1���Z���{q)Q
�Sq��Ǔg�ǽ�Dڅ&d;`�Bǫ}�U���M!ڴXHR55��,O�� �l��r������э�`-�t���[Yҙ�o�����qӛ�!xM^$�"��\��C�������PNK��/��6ʧ��q|ù#SЌ
�镼f�nVN�}��e&�7_��s��.�H�G�FC�)m�t�����ϱ��W��L�$�B�����Y=�CyY%�U�d6l�cʖQ{W�^�Z��L��p1�{�.�r�p��ح�L���%#��a|�5.�/&�b��c�^�-���>#ˬÝ��{�tq��a?�T���\5�@�Ǎ�0,��*�+�)����c��7����F��6�����A����s��~���?��eYI ��V��kSĤe�;�J��>`��(��ƒ�'���%��n��M4d��Jjꗡ��O�y���|rKQH�XA&F���.Fl������"؝'T8"3�m��
�o2�F������W���-��,�Ib�D���ٸb�%�:rL��?F+�f˛mh�0�e��?QpO� �Ih��b4�̻�"_|��9��+�bTZ}�M �ƃ�8LyYb�v�qBǺf�M����S�OM��4�g�ʂ�� �ߺ@���)�9$q��ʰ}�䷘��$#!'�m }C殦��`=����8v�9E1�2��?�x���=e�~׃&�@�q�Xb����2�)��[���Z�����¸�@��ծ^a������Կ�Ϥ:!��)����p���u��%tF���k�Y�)���A=��N�e�s?�$a��V���NѲ��V�pZ���tE^��B���i3��#�O?���q|�P�ī1�F�AÙ4�/�DD��ܗ��mntF���ϳRؼ����_˼d]&�y��N}�2�=�m�@S?�Je)�ao���f��A
7���I���w _�y�y;�Σ�FV�x��Z��'�=���aq�V�[$�n����B��$�`2�����B��&��͋C�[u5��A�407��Y#�Mʨ��N!S�3,�^���m͜?��G�?��
!�#���'��<T9�Xm�.C��pW��bv��,�
��bniA����nqHי���f҄=?�X��ڋ׃ً�Y�U4���^&�	�W����l32��;_�$|����t�� �S��j�%�x�_��ɍ��3.=��a[�)��h��/��tEJ��7�x����O:v=3�I�I&m
q��;��|�&��3�%M�'���m��ˤQh���­��5̍��Tr|���=��:�"��"�i�����F��<,ϡ�w5�t@��Fo�_�96y���hX���C��:% e�L���p�i�#XF��n���bb�α�r�=�.��W�fI ŤC0'+N��3��QkxhЃ<zV騣L��dwck6k�x�F"ra�(_��|=�w#�{G���Qg\ʊ�p&42�5a�t��!a�5"h˞��4A���Y�?$��W�פ��\ƣ��	���M�h�P߂/�͂g�c����_�صwtB���p3��
]/�^E��������'*M;V�*������ ~֯�1{m��y�˙Aн��;�y`�� \�W�}nʬm�7�S���x	�w�~���<4<+@I�3E\��ac��8������X=�hA�q�_��@�賅|���*�1�WW,}��i�&�����J!�96�<��j��Μ���R���U�ʙ��e���}5��;�?*����T�q��	�R��&tF]{�ОF( ���)Xm>�>�Q��RY�P�Ta៊�鎂$L���9^t��s�?�I�����Ӑ6�ju�*cʋ�V=���<0mP�}>��6�=3}����a�� 3�`g�LQ*��B:��.)��SRq>��!�|L�,��n��U`��E�F�f�a�|�W%
y!�/�U���qe�*�*P�'Y����ZR��[=�RɴO�ʴE����!s����]$�N���ɦ]]Wp�����)7p�\LR�AYXq��=J��$b�o$�����Ї�Gf��w*Ә6/����=lNJ�!�9��\[���+�;V͎�3E@?�/y� ��r�r�N����#t�J�O����}�tvE�K����5]���Ep5���@�v�O�&x�X�l���F����tq��3#t�l���Q��oɤx�x�7�xʁ��RU���bT������@ʌ^_\q66ER�]�x�摚1��ɴ�P��Q'����w�_�.�s�<9*��јR���lS-5l]qҒ� "|�1����g���廜��r�I�'3S���ɝ
YPNxk�ŷ��˼�.�@N�����-���������zH�o���U1MW3ޥk���N�$�[@�6`�P!J92c&�ÂAR��g.�>Z�j���&tx ��=���aOVF(��������G�b� ����Ǚ�����I�K-��s�3&p�aA�����������H(D+@��J�5ҕ�Z�]��Z��c��Ft��|#q7�����
jmު�{�QJw<Sd��"����HG�>���d|����;�#�od���!t���%w��A���ЫV�dx���i�5�n$� yK��r=ʇJ�	�r��D[4bh����?�z��~�����0�w��8�B��HC����y��)�l:+v�vB̫�;�pQH�ݴ���k)`љV� !Hz(U2A��5yq��^1l��L�L�ƻW܇�2��t��Rp��O�os��	f����rvl䜃�m�s��uŎ�\��N�����4�}�=cAi^�	�A��m�A앱�����4���qBr�����07F=��]1��X./��҂|���O�gQ|�t����t��o|^�!�(�R�is����[9ڈb^�NQC��k�g��V���jҺ)���'�Iի�
j�&�������!���Y��0�����Z��8�����HlA$2����t�n���懀_'����O	Y{>�jzx�.�JŠ�E��#�[Lag���2�������{>^s�}��,}9�++��hn�sa��O��IUC����^�r��X':�9���{�l����婔%"xEd\�gFI}��*������_�4���K������O�|B/Ҿ�����m�yDRw�=����W��D�QX� *���7�w��1�nr�z�P2�@
����.9�X�MS�!w@��N�2�?����^�PQ�4^)(UfiU9��D�r��h��ɛ3���
����=E�c�P���0m��� Y���}��)��Iޔܣ���Fq�g���}��ּ�^�>y�1~�"u�,��誮��.i��dac��bʻ3*���9��ɢ ��@�G:.zqB�n�+%}﩯��Q�_���pmD��k���M���[`D��Ż��7����8u.��1�F}"�n5�p����_�������	��"�_J�#�N�p��H���;8�.���@t�|�=i$I����P7>P�P}����d��}�t\+��3_�h�<̧����G�숞uϐTh�+=C�s^���Lj1i��Wnhk�q?s6Nt	�!�W�tD{��C}D��k����ľ����,��Ԟȝ�w�c$ps9�ޣ�M�|�x��q�[w���$e��y�ײr���g�?$�(�y.I�tx�S��-\�a����_�<<.� g�����%z= �'��u\��%�|��&��/z^��36^���k��s�c�R��`�l�h�� ��(SI�Y`,��Hk�6�Z�TK�54H�^�ˌ���D鰫�Uw��:�a���Xg�}~ؑb�����^��c�p	_$�I5�^#�ɤ��;/1n
��'�9\��!���|�H)�S ���M������^��y Z�T�kY4;"ӡ+�+Pf
���}���|��+G-�y�X���_#6�yC�HZ���V/̲Q`c@�����:���C���J���V�ͅRl������'�{'�_��t����7Z|��7����bx��l�<�,�։H3nL_s�ŋۭ/Q�{H��Yk��\-i仪�ǧS��R��%:ܭ -��6����Q����0 F�+%���Zaic�����P���@$R����d
WR�])�&�5����BoO����x�A����@ݜJ��f��νI�X�� o$�D3wr`:���"���.����z�`��ˡ
���~������ِ�ѽ�'��Z).��\T$�`�V{>�X����|�?K��,�P�&G<B�
�6ۦn���Cඦw<�AT�%�ަ]?P�e���������0��
�n��r��A��2/���(P0n!�\|�i⢰��[�Q��e<�om�
���f���avEh1��e�,h�b<V�)�UѴ��X:�s0�|�m�9�w@0�va�m2�"�57�ן����
����[ƛ� �2�ٯo|>z��$۩Æ< ��ԧ_>Rb"�:�o��9fdo�Fq.ёwּd�(?�����9�k/�<�O!�A�"�G���n�K,���봔�G��� D�Za?U�jj�A`=�$<����S���2(�(l`������9[P��Kh)*�F��E3�7�|̥]������[�a��w�#4��=�Q��ɺ͆�L�E��хd[䔁��D����Oҹjŵ�g���1��mgfJ��'=��ź�rl%\8��3ʷ�܏��^�Wgr�3�X�w�e�YY���i��X�??��!�b�r-�`�fɊ_��7)�iUP����)lM��X�_nB��a]����Z�
^���І�[҄��#�\��j$�$�.��9�D�F���F�Lͮ��y���qT�bD������pB��6R:sq]�Mi���e�À1������qS��W��xh*��c0C�����Eqȶt���5�൜2�_!"6�B���NWՉe�@��5�����*>q&h��n9�N��$�Z$�TE����%��寏�n2(I�!�A��1�[���K�N��1�"X�F$9<Hm,*�T�x��e����~\CC�L�]{�g���I@WG���$���B׆t�^J*��=�"�柃ul�Ϧ�5١u��?�ʜ��<���X��!��h�*��_KJ�=�!�7;�Gcw���{����)�l�G��s�"�i����y��d`�|���]O~�B|��s��<�{~�o9�͂͞��XG[W ȯsƊĩ=��ZKg�/)�K�=�unx�����S��� �γ��&r��L�1�2�^�"��Aw��#S� Ļ$�ž��z.�~��}��V���t�	y�o,�AsM^X��Π������Q�T�*�eA�P��)m�)�g�ӜN��1oj�Fa�&p�y�r�ĵ�D�4�!�����7b�2x��}�q%���迹�7�a��7)�z��&$�æ ^UYf��h���
�Oĥ]��6��NN�ŠCD

�}m�B��1.�o����=n���V�!d�n��mO�N�>v>}�)�<2���)�ڃK0�q(�C8�S%�X���q�'���J�i|G��>���-!�hf{�9V���«�%�ok�����+v��.o<Mα����yԌZ:�q �z��\nOK��]�b��	�*�����_�l��fn���b�Q���Z%�{� ��A�S���Ԓ�vv�\c@!�Jܭ_uh�2(Ȳ^u� ��9��@dƪ�Ž�,V����]rl�q|��ͷ�0�Ia��6Y�7A-�4e�
��4�!���*
�8� 8�����%�/��������1ja���W�r ��a����	�}�I�PF 5�^�,�s�iH`��K,��q�$�'�Ǘg���j�o��*DP��C*�t���!E���u��n����w]m�V.��m�s���ȕ�lY�����	����$(���䟂o` X�o�QF�Aϊ����������/���y�����!KXX���)�?���� D�,64��t��
���>��i�T���綨zĬ����I��`S'�S��X�r! ��Y7nL%:��WԀ��qԸWͰ��y���^Me��k��1b�>�����j�%>��Ӻ�/�d�a�" �p<�|N⺓�3R�����w.u���=��`AbI=.��x��df��i�Q��v���2hB_C�j �"Ƃ�1gux�o�x�H��)rz{��p�aMd_�Ϥ>X��C�E�����|H�v����.��Å'#�Lɽ񊢳��?ޛY���1dVPK+T�Ϻҵx���M.e����8Ȉ���[(41&oA�;��w��a.V��Wl�G����m=�f,��:&��1X��B�rm;d�����Pj8�^8|�5�m�y�b�����U��~���R�������%^3���;V0�����M�1�	i�P�P��?0� 5ҏ�����3q��2��4�fi��/:��������Y
���DA0����(��腬�۳U�h��o���+8ǵu�-�nUj��i��.���eJ�cZ�E�QUP��ω�`�X�T ��ATd63��Y�^�d]s6�8]eq�?�����p��E�yO����|��r{�w�����'����0��g�B%Is����G��4	A�ԃ3�]����n��+���I'�p<�G��N�����5��p�|�ucf��P�%+<K~pY�V$\w���Sj������CM�f�ǐ�6>��l�����	�cH�U�)u�\{j�U��R��e~t	
.~�����]+�Q��J8+����_���}������C��@6ŀZ�`�2�'�����*㤹j���YG��D��!�pY{?�6Q����V�.I���t���<���c��*�c��( �"�)��Ez����`M���-����F��n�՚�f�11���%��ʾ��0��W��P >��f�]�v� �� bQ!|�FK��C$��G�+ZP��b�v�?j�X��4���>f�N�%�E�0N��dX[�� S�Y8��\6 f>����8&�W[�A0�[�}��s~qr�	F�z� ���4&�Q��N�*\�G��g4zh�f�E9%@�����
�r��?�:��gv�2�<�eo��N��}w\��_�ΊӴA�W�W�yKUA� Y��o#@vؕ�Z ޷�_��X����7��[�9�Ջ�v�=ǔ��{-�a�:r�D(Uz����;BLY��~â�����֪q���~��+�I��m�*�f;�d�>
79ZO�vџ��Iw}�!�����ό/�M�.��-�o�V��(
����<Q��گj��~��m�Y;�@\^�����mGT� ȀCIC�G��o��dB�=��	p0`�4ß���G��`���� `���YLad��G��τM��P�4���58͜�K�%z���"����{͆��?��y%��ϭ������L��ќ��<�z����,�U���<|l{