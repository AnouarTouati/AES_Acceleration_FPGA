��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pٌ9=��	�[L�⏥2��֕���z�Q1�A�����p�
�D�2��rͻ12�mo�Xa�{�c 9�������0��]��R҈N=����cM��H�-v�ބ��uA�k���=Qߋ+e$FY
�	HZ��9liolNCcaty{#Q�?�|����� >VRw:nR����P瞮 o�K�3)怒�6n"��{�ͩL�{_���I�Jf�9�\�m���HLH�f���w�t��fhq#�~��F��m&�%[��<w��VS�#�3����}��j�z���.5G��#�z�Em�MXnJF���3|!����ʼ+��`�da�3���;^��ĠJ�w|��D��Ҙ���-��Q��9�Q�z�����,j�!��]{q|�x����qS薿���,�%2}��	�#vF|s;L�"HF�e�x홿Y�.���#� ���W��1Lte��+0q�#jC����+��!#ҭ����%h��iwu���3����?����|a�ݐJ��R&L5�$�ɿ�֒�Y�Ę9P�WKU�qb5#D51ȰdvŶA3�S�"�a�!�M�K�ëV���4��лz"at�n�\���}wm�h��9�qO?k
���e���i*&��!H������`�Ci�Ǉ�$���,�jp�8���w,��V���/h�|W�x2�E:�zK��k_�����#ͧ+�U��o��}Sq�����O�+4c ͌�͈��%2�v���������77f^�嗘����'/�1�O�h~�L�����Q"��KtJ�H�F�t�M��.i�6���zHP�z=���Tu�*;z�$n��=z2z��ő(�;��Ǌ�=�u�o���h�R��=o�r�4~$� #iH܌o/F��$鼎���{/����k�β��mÊ������7C�w�!�8*l��T���ա@���H0�[�W#=��JwQx����c�P���F��;��2W�vR2�����*����&�0�����LcJ>��Î}�V���ktn�j�"�T�a�Ub3��c�&)�X��z!�k����k/	ʋ�tL��1N���'���XX}r���6XNH�RR�?#}p;�MO:��Ox$v�Y� ����K����&��.mC;��D�؈�����.��Pax��1��2���{��.-^�W��G��z���O�b�M�< ���->?N������#�[pk��^�Ֆ�#��u���
g${�ˤ�B���g�����.�
�ޓ�o�/,������".;��e����0�XU���J���/��г��p?�٬Ecӗ���I�K�?��6��_Ew����ֵ���֗���Rc����f6�;�P;P�#�t�wg�\� I�c�C��8g���c#����_�!J�R�0�&~����(�}\��W}-��s����W^~|���W����Ɗ�R�R��p4J��xN�=d�"L�bq��}�!A��cZ�ʿ�^h;L�<Ŋ����l-����M��2�.���2'+#�\�هw2��=0����&y����i��-�R�W@����?$�2Cb+�VoIɆ�f2�m���� ���_��B�d�8JI� N���4�:T�՛aVx���v�І�o���Y��g�:Y��j��]�B�o��t6SG S�oG�7�\i!M�L'������4�r{�V��z�P�=�7B�����fl���@��'�y�L�����5Ax�3�P=E+��EN�i�w�����c��x %� �]��w1�!|���W��|j�xv+Q[AԸ&��ߡ��CI��eO�C M.�Aܽ��(S���hV�_?6�l�r���
�^~�!�b���	]1��2rK,d��~�U��G�J����i�=6���X:a2{Pr�[�zi�b&D������ȫ'D |ӻlۮ|���_'����ʖȣ�� `�.*� �8*<��|x��z�ͷ������)琢��B�
��];�	���P�m�s����!y��5b��?53�\c��@��{)��[����è���Xq>���@W�T'�cg��.|���9�w�uh��<�#���˳'�y*��qB����u싗r$�M�k|�j����>6�a��x	q^7NсZ�y�����\R,�@eŰz[^r GvE�o��+?[$^�����`����7���)���&G�!�<�e���M1ݾ�0�R"#1��<�������v����X�[�F�g�2���2��c��J�6/�jM�a�&乔���WH�)��K_��d�ft��(��wP�.���S86OBډVx�Ga���R��޸�p	^�ja!��N�a!�o�m�<dz�SZLm6���R>:���撟�%��R���D�e��/�!)�5=3�K������Z���㖚Tw��2��^9&���9xs�����\n���+xN�={Ƿ���k�+���sY�7���M��C��f0VR���Z���Îh=��a=��;�'���)�����(}ʓ�9�hdh=&�����E��<��{���~�ϲ6�%#ͷȖ5vomy�.2p���D����[�<(J�0@(B��%��	�ao��ќ���k��w��vnt?n�{�v��R�PUt�[}��	-��I���'�4j�)���v=B�O����x�]�[��\9X;s�ՇU�-h��Z��b'���)��M:�l_#m���oykIX���>YW.����Ҷ@(sir�f+���W=����Bh^�SW%�mqx�$��P�{lK�W�r zkw����pXa��e3x0魅��]x>��w�
I)s.�ƬO����
!i:�Z�������wGB�j�����#�G߉"�8�|<c;Am�����{��)DW�Qm�tL� �Q�a���jj $�n�+E��Uʧ+����6::I�#I ���q\�p������EC��d��~��V��A+̺�Α�"Y�]>�����m�{/" ��Cob���n2�'"0&�&�����r#��UzR }��rb����o����^�!�f]*�X�;(�]���Y���t��y��g&����V�R��s��\�T]]�z�w�_�o�zG��v���lp�S�a��x��=fA�Bx2�8J�3�l*��5����;��?���	?��C�Q4b�ס��,9����P��\���@�Z�����r.z�b�cj�V#{�f�[��^�E �(�P���>ƻWX(�I�D s��^��6aR �ؐm-�u&|�\zi�19ْ��V�X�������ɺ4ݱ .-c��K �E5�mEl%��FT;B����7�n���`�)��A�+�`ts��*/&F�8������;X�pB)	�~���{8N���%�i/�YZmz�e1F�� �,�=W�i�8o�P�.��o�)@��ZBf�c	C �w}R`�p4�j�츃��-��v"p����כ�%�����	�mhHZ�QZ�EY�A��+��~���2��� �u �CB�DQ#��?�aD���M�_�!�	;x�۲�BH����"�;:�����0�����-d�����(^'�/�`O�N"0{/Y����[%u���X��������8���@F��-�ߢ��cHP:��Q��D�X�����O��0�p�;X��x�Iu��IzBv:;w�x����4��O2�d��{�٨=��S�a�)@OΏ,e0<z��lZ��s����!�N3�2��WS�d���"���HX4*M���כ�g�g�����%�U�3�#��>��V ``.:�t��D����:�aS�N��Y_RTx����7+P0�IK"��~�B�:�p���T�2��1Z�ۊ,*��eC�t��j��٬�5"��e5��9!`�WH[�� 5'2*UK7�º��G���®HR�zL^��T��/a�1�yUI��⍻�<b�1��'��ĥt*�0!��s6v��~5�h�7�����ձ�{*J�^1�џ��92�?�~�R��EMO�yˮv3N�8��[�-�]s�!��]ƶ�70�l+�XP�ո�����.{��(E~�7rԣw# U���~��i�Vs�}%}��Q�3_�����Ć���Wx�
�+�GB`��M?xSB©z����,�����#\|}#�Y����xD�,&�"]�	�� V9,��0t�Į�&�8�Jh�zt�4pZ��YKo��#ܤ�=x^�Q��!�݅�t�N�\H&(Ky�	u�M$)�y��q�ǧ)��#W�^�_IrѰ�g���$��v܋K�וSs��ZDX���BO���3��ꜥ�G�g~ps�:ܚA���v�VqRy���[��5�<���6�[;vB��J�R>DXAPk����#��&��EZ��4�C��e;K�]C!c�89�����f J݇&0-�s�����0����W �$��\I�����_.�$�l�N^�=�7w��S{w��r\����
�+d2eB�6v V�|��g�����$8�/��N� *85����2���\�-]Yn��9���� ��{�EtR�-��u��L��3{��u����-�J��XroxA��A�冉nn����{����������l�`v����]DRx
ՙ��
֕���F`�e�����{���h�B:��7��O��(�n������U�SH�t�D�'�k��:�J�����/��O�W	pT���\Bh4��2eL,q�~�/gF*��f�]Wt�-���Ee�~u�zjb���r>�R���{tβJ�P����1ABh�m��?(N*�㬣�Z�4s��p�@i�NX�rvx�����$��v̷qghf� ]z|����h�ыI��n�@1�v��"h��%�)O ���+I(Y��׀��a��`X5g�-��Y_�=ax�b�u�'74i9!����sܦ2R?�|�����b���BC���l��v���m����2�&(3m��y���}ʃ����9ad�l�w�P�w�Ű��E�cH,y~ofB`��P:�������� '�Nw�<:^iz�$��W�p�~����a�Ǒ����[
"M�ᾉE뜬����ֽ}�+ ��RJ�Lt��0�~�p�����kN_��8�o����51P�&�Y��&4��fS��� U<���!{GCو�}�)�N�$�GX��yR�Si��搻�g�?�sPe��sh�\��V��hd�U���*2ט�pԸy��#QsRM�<�(����@W�SUJgh�J������Z��-쉣
�t,�~�Yy�6"��>��䀜0��v�C�DY�0X\<��5�W�&���6E��!���Nʹ���8]U'_�����!��Z�֥w�+cm��]ב�{1��{�{��;�7d��ߵ[Cma@m�3 �8b�B��k�h�����4U���c��y��j���plh���>O��͛|gkB>_�l����gU�` F��y�����2�ف��.Ș�5@�S`�0�%i� �9���nD�mg"`�4u6�D�������w�>6����Ӟú�e�$��=��j��Jo�����˘[?rQ��k��:��Rk ������|�����ݷ_7��-��b�O�b�G�Ue�������B�!��	~(J�O�w�awa�������ނ��g�5
���^��h�J��;�F�o���qir{%��=�k6@��ѲG�b���o��;�m�Ѳ����p
�9L?=Z5�[�̓�������c�@!��|�ά%{������{�9���M���c�<TM�-^���?N�����k���7/�O�gSJ��fp����d��qzd�՛n�F'�pa8Y48��8����e���O�8��4�:�h#�Dj�U�������n���E���+Ƶ�V�WR�+Q�:�P8�f� �����b�䅑{tǭ	ĳ�G� C��d�����0� %o���[�p֥(=�y�bc� ����Q��M�GkxSv�Z|�o�&u�8�:�UW�N1�W�q:���˗	�fM��^J@��C�s����-uΤ+�'��y�IN_�ߓ0(GsR87A�F#��:����Z�;��<"c>%|d�@�U��M������ւ�yµ�Ψ�.]`���;>��w^E������!#C%@�2Rň�����dm��Y=�q"�.����D����%��-�.���7���/���؎w�hw�n��2r8�Θ+O�$|��O��E�!Ą'(aƈ��4o4����]ܵ����	���7I�UA���r�ıv��v�C�� 
�h�L!vс��?.��&��<�K�E�r�ްl���S� �g�',���꿗��>�]��?�ƴ�u��#��BAc�������=q��r�)l�C�Iv�qM��'�+�Q��޶M�;k��#Sf�gtU�tUtAT�,ܤY���}����[�RJ}s	�*�F;O����\��t�*����l�4��]W�\�_~^ ����g�1M@Y���� \ɋ<�}®J�!��7�g�Tf(xv��?<�J�ݯ�N�*�Ƶ�o��Y��lV��o��wp��5������bW����H���X#2�$�����A!:�� ,���z�P�IEW���	p6��Z������¨�;�@2���+���J��ˠ�~ �M�c�733�M�X-�b��Q�_$���2��ۗ5�b@�g[)ߤ{�\m�pj��mwn��+������q�LACc�y�1C$6�\�lkzL��.�>?�a������.�u �k��gQ��`>�X�H�i���mN�j"
��ӏY@�����O�Y��({�JY�9]�ըMN�K*��������X��Yإ�W�����J�N�y�@|	+fZ���{V,
�E]V�y�eC�4�1rwPX�TER
��b*���\�5jh����y�^d���31[8R�����3z�!���"�=��]~�H�/���#;������r������ߤ$n�zT>��:�{ϑ�J����^�:�A%�Ŧ"��\�S���z��륝��,k���?%�7��K�AJfM8j�W#l7{�i /IBzM�a��H;s��t
��ێ��7x��x�D'h��5O��)�XFg���N�n�lT��~�x�Tn�:Ӈurߩ.���5 �).��� L�D�&z�'>���!���Gp�/geǶ��� 3F�W�����^�9���K�`�1�����n���D��;w�=�^!���I;�Qz�FJW���u%Ͳ�]�qV�]�)��&��Xg��Bo6����a V�L�Za�L�����;źri�������-� "�n���	G����<��$��gb���2�#"�����/�Ok*���i�X���lq������E����{-5@l0&��ac�7#V�s%�ON?؏d�,
�|�0�K�L���r�{k��(�|uS5��[�9I;mf�a"�w�E(���f��>[9n���DR ��0���w�5}�(�9*w�L`X:�&"�1H$���by����?a���H�qnݹ����IQ��͎4Y��ߘ}��Ь/FU�]k��p�:�ՠ�@�)E������G�6B$���A�oJ���Dв�eW���?�&�i���r�&�K�ا�ƕ;���)�{��2ێ�E�
��mtվ��m�l�q�}�kЕ��l����vl׻]�	VH�=��z���;`ts$@��T�غ��5!����� q l�&�/(F�a����i�6�U'e=:@�7齗ؐHmx������|��+D��[��Twd�<o�v�[|�IN6�ѩ5� ��&�`�-˃�]}���ao�nd�w�����U�a�G��އ�V���^�)��f�i����l�Ck^���ߩ�N\,Q�W�����L��(����g&Ņ��BP5д����!ތ��6�rBes*f���zjB����g���$�t?��[I���-,d^L������HF3#��;K���g?3a�vw0��-3�}m����%2����T�sK��;�g���!x�rKF�2��\Ŧ���&���^?��$�,�M�g5?O����0��p-��V�9����p�:��H��k��TY���J��/��<�bݻ���<�B�\tF��;L����__��L��ø�s4���B
�d��������T�ʶ����oIg���Ԇ�=��{м��F2���B}o�0�y�ev��	���e�u"l܎��k� ;��{�ՈM���B���~��5��Zhe�� <��b��a������A�x���>ơ5��M>�=M=��ǅ
�z���毚�A���]V�yi�@� ���DP�b�O:/iE�H�A>d����Yd��*�"�B��xPe~ (3�7��a˅LTJ�# v�"L�,���"�@I�
�N���)c>s���#~eB���J�Q�ug_*��-�<�����iҗ#[SAܯfN�R�����>���o��i|I��W�	������WC�9� 	L�U'�����jW���<~`���8��"z�M����c4�m����:��fP���.� �
����h��n)Dv? �-��&���KO�"ޤ�c;��$:��9:�?X������>�<{�V�X���B��h�e�i�Tv�6V����M���v���|��r����#�čz��^��H�w�5������ѯ�9៊���&����Tb=�,���/�����;�d�� �}�ϋ�h��\��V(��� 5�z��x��w��!�"������(��wi�a��5���pep�K6����bt�̛wNF�M�<�QOa��[(�b1�.��Kg���}4��s1�cgC:�u�:.@m����|��Đ��H����+&��E��q)�Cs�JAjG�����>R'� 5�h,�93�7��6��"d����9?a��G�l�G.FT������	
�
�7rE2i��)"W��L��Qn�$|�j`����v�bAx��~�%ǄP���Z��Ͷ\�v��:��9w"�CׯR�u|�c>�=j�9r��J��<��-���~`�e�����r4�3!z�l [���ί�L� �=�A=��D�8q���7��.�OT;�+�/�äsL�+Q�k�w$� ���6>()IN4.�D������,�SJ!̤bȠ$��k��t#ʦ���y��c�2k�`8��������N��m��8�"��6��6{�xf�8����cVl7G����O�3qt! W��2�7�p���Ը�`��i6��j�Ffɲ�_bR�L����8�����;&��!|�]D
�2���)oB$g���A�h��A�\.��r�܋��o_��L��Gzp�Zb���ܼ9���IsW���P�5_j������G*W�Lp7�Q�ӕ��)������ʨ��"���Y)�%ʤ�>�Q�=}��7�	`��?��h�Ĭ�e2��j;vT~��M�(Z=�)������\۟V�=-tϊՓ�Fr=�̷�)��#J��	e��+U��Q�Fj�桏н�^<����ԋ��]���6�>��r�<�����#lq�La��v��>yD=kO�$�-�y���v��m�j�܀�%X��L��[��6�ݦ���C{O�%�n�PS??�۪�ܐE�|�{��,�����Դ����Q�79��E��&��h#JC��Y��tr��)��F��
�)Y�mm�a���O^��{���Q�^��v�f	r-%�{��8�X�<]�+������ۗ{��htv�<?ZHtk�t"��C�iEM�;�^������QV'�F��A��U�C�w
H�{�Eߛ���02�����K�Pq��41�c�]��^N똑���p�ݘ/����ٌ��˫ӗ��o$&�� G�����~g�z�W�k���$~q~6�#ʗ9lK����:8C��.��v�wpJ���t?��m�����8a�C��O��łK����
�P���-̵(+�(�K7��#]k��:_��er��%��
ƭ3 m��hY�7�G�Ci Awk��/�딥^��K����:	SݶJ;.�m��@H��#ù���(�Y��1h�J(?�~�s�m��@P=����v���ҚJ� ���HoR�.��T�8�j��w���� �|j����ɴ�E��V�C�l���i�6�O���w<
�ޟa�TJ4�-ܦh�I�Z�n�M��V8�<6zTm@�X.^�D�݂7r�4(��L��d��yi0��-�90GI7n0��6Mb�{4hF1ץ�g�>N����s��̨�,_�$`T�2����Q~ƭ[��j��p4�Q��&��ޚwO�&"����� ꆷIJ*����
?@��]R���gq���c��!��%B�j�bhЊ��8�	��{u!�aR�7��k���YE@�)��-hb eۛ��(�f�vk�i��ղ���f�r'_W!\g��+���$�����>v.���>��f�s��HM=�����D("��������[��]�qd���S�G�(�Co=���b�A�t����Ⱦ5��ϖ�J�3�t���?�ڒ����*Ux��b�3!�nH02���o=����GK�KG�	�~YN��4m�p�1��r��s�]�f�H����@d"m:�$����<_4���g�\8�d<Y���2G;��_+Μ��&��r6�F�F(��dRnh��4QC����bJ֨�� �ߣm�������OBOE/�>N�:�L��Jқ�"zB�0\�7�Q�_<��MF)�� .f
!<���Q�I��T�HT���N��f&;����|�X��M2�Z��q�&�r!�e���q؆{	c�hE9�/�ZxJ���3E:睎�HЖc��XK
i���'&^���?:�Y6J�ҟ�n�P3��77rIHt8I߄+hר�7l"㾉���Op�3��H��g9���1-(:c`t���A\\>=hptn,{E@j_!uj!�1N��CkEl��x:��TH2|�M���v��U� Vrb
��v�����MP '�XhQ�k�L����q]��p��6Թ�~vA���ǐT<u�	������.�S%�#w%Ŝ|��v�ϼ�F�du��U"G��
0z�<[W�_tR�N�b@>��?=�5��d'�Ϳaq�@���q5Z��� q��n��Iݺ�9�����4a����5Lp=&Pfde�M���aߡ�/����&9,�mܱ"�n£������n-��V3���>j�����
�m�:d��	�ޭ^-����`H���c����flʐoߊ,�2��ZE���{]Hh4�OJ�R��1���7�.r�|w8t5o����t��@vľdS&G�k�.JQ�ϖѵ:��g:!c4�3�IfB���#3wjtw:8=�[̣���v�ͩS�f�.�\8g��x����[�Y[����śǼ�
s�Rt��؜�coeXc]���/:?�K1׳��BIG|�
�����fKF�ީ�k<�v�s�O�r��տ��a�� Z�$��G����	�˃{�-����V����QI�.c������} U����.�U �I���>�����H�2������R�z�w
Г	�O%��L.��0q��ܚ�{�s��q8�V3];�ӌ��q5�h�J��l,<0��U����±��X�t"T�F7�e���z�Ǆߕ������1#��{Å���8��s�m��{��Ў�U0�H�
����R�°�6��Z�Q���Sp�&3�F*�����́R�(B,��'�D{��xI8 ������c�s�P�X�j)] @ӡ��˧����AŘ~\�b��6��8���X�/��x \�v��1J�XD0�,����@���}�{���so�p���/�j��e{V��-�,�77��-�ו�����t )qz�w�����p�gND �̽�TU�{Qt��/�ٌdX�1nc�:(k�C���l�2&��f�`�[��9XR��P�u��E$VDy7����x9�;ts��%>d\������l�����I?�@��(���F�w��]���N�h�A|-�梥I��(�o�P��[3�mr��e�΃��_�ԟ�|��{�����;����}-�D�؆��G?���pie���)������G��o��Ђ�u
Dm�ڙO� �	�R+V�a��9��H
�F�_/��U�Ȋ�_=Lu�Q��\w=�N�����"���[ヒh�Y�'q̍j���{k�q<8�΄��௭�0o�?�r�|%�x1��єl�6|0y۪b[�����5�D���ƃJ<�}1^�P0���_g[���Ca�C0*ˢ�e�����-���T��R�8NQ��L:=X%��T�b�cI�O��h>uӲY��>��h���qM��U)s�'{���PH��	��>`O�:�5����c�4�~�O?T�y\)��엚|خ"`ҤcO$=�[��6c�ǭ�Z-�X��O������Ė��R��.�"մlz�$??/:�}�U�����Y��{uX�B$#s�9B��ǂ�w�hB�j��Ω��M]Z�i]�z&.�#3��\�ˌ����Cl �N�)`-�T�o�gW�n��c	���o?~@
�X*�y^bi/�:���	��M2I3y�9���7��k�D;:��D� C�Qd�e�:XsX��=|둩�qU6��Y�_�f4x��$�a@�����.@.z��%v`d���^�@�����b�Nֲ��惔�O���!Mu�V[P�#��srf�&��)�0�W�|�M��?!/b+%p+�������C	���Ԟ�X�K1�д��&�uD����H�� \w=��+䆴K'����0���y�㖨�O��T�-YyTU�Xl�F�Q�f�#��]�v/��$������~\�� ��(R!�}���^C?�Ȑ������5}BXA$O��u�QZ#^�vz��_jՊ��|"�]x��S�Ȫ�����-c���uGĽ�Ρ�/Ź����A6�'6��V�R�B]��0<hw"�p��v�{�w��%���0smHN�.wFtIĳ%i�<t�"\��8gT�f�ӑ}��r8��sAtIn=c܃�^z�d��c�DD�V4O����u\��HU�u�u7	�N�l��3�����rlr8� h���s{X &��h0�4�_� ���k3�:�fk,�Z�# CT:2N9n��v�/YH�Bp�$h8��z��.
H�м*�\��|@f�TG3l���[<�Es�,�+GM?5։3~W<]Dj��/�|z
�
�s�Y��b�	@��6�~g>t�}����u�l9rh)C���[��S����*k$�תw�B;̕Q(HSE�n�(�{��i�5r2��Z�q�d�m-�6�	��e�E��t��s"pj�X� A�jH�Ap��l��Bb��[R�s�	�	](����,L�.����	�mB��'+h�v�,�@m.-Rs
P=|o�Nt�)���t
~���tP�����瓣�&�~��156S��xm ߧZ�^}�.�va`�쬍n�x�d�<rAX�;T���Z�C]_K����F�X��v��.��6��,��R(E����K"G�J�;�B���5�����lE����f�z�λ���Bj�%����bM�Rٓl��~��vW`��$�]&����Rxu^��h�`�	f�0�0luzP�'�3��!ZC��T+�ώW��K$�+�v.AX0���ѐ#/'�&��!M�U�d�h%���<�ER"�3��	c�õ�;I�w0[�J�����M�imݘ�%��`rd�4fvn}$�h%�
49����=f�2�D�n	o"�-&ǀC��DҺ��|p�ϒ��/����Kx^y.Ǖ�A�. C�J]ʦv/Qǂ�@�ΒA�t4�V���� m���dx��:rݧ��0�[�^d���Ib�����0a���ǣF�h������#�`q3w.[�=�MZN����H	X&���խ���)U�T�Oa�N�F�)�E"�G��i�Э�*o��b���yB6����"����Zq�nHi���ɇJ ��'9��	�W�
Q8�,^�PU+<� ���b�3��!��F+�z�����u�W|}↑��T�E�������eF�r����6'p��ӵꞺ�9��a}�[��0<:*�/�ETW�e27IIn�/�+�G+M%dBhp���$:��J��T{��z�vT�:�~���m����	A@A�\��D8����n����S��҆r�WP���m��.�k ����(����y��jE�i�BY�1�xp\�1[9��+�S��O�j��8z�fS0�u���<�����9',�ȹ;c<5H�������K갉�c<�Q�z��-���n���R��<P/Z9|�����]^!�iu�\|Y����/6I�_�^.ò�l��X7>x�b{��,"�|c���#?��oɷJ�dˀ@�o��2���;^�'�g�����82\��"K�Q�mL̃^��k�q�����0/�i\)��cN��
�YW;�z�oW]�N�v�sj��P���3	���'������e�=L��훶-�η�p���p�DI@_ĉ�FOo^���}��؃	,�?L>9��,���?��]=�!��ϴ�Y��籛�"���^�����S-wtt�st�X�R�g��g|X�Lx.o�r�*8�G����$���[��{Su���%Cop,׾�9�������L��;܎�Z0u���6v�+�%�57;���y5lY8'3lW��^�1���ƚ��lI�~��W�q�S�.�XJ�oåY��I�~���4w�*ߦ>߹����"�h?7�Q�����zd����g	���$9=�%�e�OH2Y����l߅�0�����jQF�H��R�y��f�n��K�)�Ӂ0���f��l������C�q��0Yx�9�����,�����g���Q�z|����,Zs֣���j%�$m����K>���Z��A����MfQ����_-�3�/y��Vw�T�P���T�: ��]�[Q{�}�H��Mw������,�"؃�
��/���Ceq���+�o��˫dB�dpσmVu��Gl�sf��k
�
z��u,}Ͻ��>_�k�k�l5Pǭ°z���?���3��S��hxl<�#�<�dO���I�Ա��^���b�(�uF~b�@�w!I� �9�S���4}��],sg�Bb	�8&��Md��,�H���#HW���&n��E�#���"5{g�7�9�H�!�w�Ĉk���������7���ڕ�?��f���-Ȭ̧���q���1�O{� �hq�4r�Q��آ�l�Z��K!��e�+�J�tJ��l.;�`!�򊠳�0\����J �_�=�n ���r�Z��R���|dÕ��b�h��c�$?+(�3g��
�=0�T\G%���XL�E=R0+����,1�=��6j>��;�{�zNn�P���r\IZ�,.�P��������#D��|�v&��EQDKI	LH�	��4�[R�[�� xA�g�����-a�����G�ݟ��=n�z�Nk$Gi��X#k^�)/OE�
3��`/t���A����2gO�rn�f=����~O��<��}��n=�8��B*V�.�B�%�p.yf�#Z����2o`g<r��}v�Z���$�Vۛ��h��|�8��%����	:�Ȣ����^vXنJO��*L�7�'���8��� ֹ'ǹ@��T^�4;{�-���:��5�YF��H�S��)��̼���[cN��A�7j'7��e���᧸��_}��y��n[r2m�T��8��  ���t����Ut
%�+Rk���
<���α%�pL2�'��t��`c�kR4��\�͏0v�\���z�����0��(�|c	���b�O��7"��(�/�'q�z;^��08?�Zi�Re���?���)�ǯ6&�k�����GE;ƍ�O�iW�sߠ�]mvA��N�{~��W[��4x9iBLq#�z�HGS��0[��~��|�:�8҈�R���h>���Qj�h��:b"v�3J$�f��(p�ђ�L$V��D�J��ޠ g*V%1bum�v�"SP-@��ӫ���xi/ ���d5�=�g=Fy[=ah��;�J^��{]n$`�m�)*γ1,��=�~�Hk�_"a�3/T
0;B�!�m{�I�������E�l�׿����f}��)����A�Ј�D��Φm���O����?�8���Q�Ҍ������p3)P����@Hz����Z�/�&�ݬ@�U!�b���\-���9��RQ�B�Ӈ���ǈ��B`Ӵ��j]f\��'���%�/�]�[�\Nx� �����?��C�D~�H��i;�V�6f�A��B�8�^���>�����r���~6+��oP'j����H$�oß\��Dߢ��Y�:�H_L=���Y����
�
� �XI%.�Z��æ��e��5#f�Ӷ��7U��i�G�ȫ�Ci͝����
�Mr~;�:��������M��E�i��^SZ�F<K�#�f��yZ
�i�z%��
.��>�|�"�	��f��*�$�
�e�1��p��r7'T�c̵Hs��=����̼D�Q�g#lت�2v�v��[�Y��~>�j"�����y�$)�V�Q�F�пF[���\P��,�S�;� R�+��T��ן� ����2�tK���/k�."�Re/?��N�Єo�с�����8����m�Ub+%�f�A��tdw�ԩ)7v��&��ߋׅ��L�F�
/*���P�F[J��F�6x���s����o=�|�������ߌ����U��M��Έڸ��xPLCE�]�ȻU�A�}�w<)���Ɏ;*���	�v��[�[T˲K����
5R�9�2~�u��n�-��7$�n�_G��k٥�Myx}P�.�-�����S���y6�T\J7NΞb��;��ּ��I�y5�J�~������O3Zۅ\O�'z0n*�x�_�zߐ��%�=���O��
"��h�J¤�Ig��N<��Ee:��oJn�oJ��Ⱥ�_��$,�3��+zA����"m��R��o�F.S��+�7�aH���VG�.(bG�~�O�R]����3�i������:ղ,� -��}}�ֹ�/m�B,�O��L�Xm:���/��{��}���@>�O�~�ʮ�~+X/}1�\�)=���~��>�"-�bI?x���Ϣ�Q~kV�⨚�&Պ�^,�!f��v�@��ր�o"BF�L����fämY���7`9Z�M6�H�Ls�C�@���z�	ݬ1c���(�x��������?��
��"���E�ӌ�����D�O��@�k�9B<��'B=�U0@T���Dx�zC�\�0��(%�:<��t@��$�*��f���Ҟ�_q��3>E2�(�W�f�o�N�P}�Y�<�ѯ��t �r	�K���9(,m҆���,�\*�5�AКi��Ȏ�w�>�nCCz�w�"�;�����Qe	�lj��|�5�$o��z�'��Q�PsE![����;����T��̾�B��1O�e��Vz��{��a��d[�w�I�Ŋ�6ETN@�u����A@v��)�9�J�(�܎x�E�aE�.���Ґ��U���Mt����dS܏�%������<O[�4k�Ͻ�W0j���[2�<7�4��+B��;��an\L�i��,���ǔR��}(ڌ��ˑh�Eţ6Sv�9м�����͒NXˆ�	�
�B��g���M��Z�<�Ĩ�iľ&���`��pg�e���&�;�`�-U�wj�mt�`}C��@�t��+�W��z�62/P�ퟳ��;�͏JXT���qA,��m�xX�\�H�������r:(RSA�~�lC����+�f���F�!J����8����<�l���~�@� ��33^[�haAN[��.Pr���G�ݥi,��Ǹݙ���] }U��mF7�m�{f�;?~�ȨL���<�N�R��,�t���������tV-�������}���L6��ִKޤ��4Ɲ�x�Z�-��ݼ3�X���j�%�M�_���4�Y����*b��F��'����-8���"��r��PO�f_7��ɾվ�V��)�ڦ��h+#�N�9Dh�>W�(��&�?�S`��#z�����)��-�*�O=��`�"E�����26ټ�e������(���U�s�1�휘�A~:HWZ�/?"!����ѥ|�p��M�D�h1Z�V�ϒd#���$�<2��u(5J���uw���rQ� "X��/�I�l�-��6�Wy����8�]g�Z�Õ.?qími'b���|3����j�=M�Q�Լa���D�I1�̆�6��S^�*x�^0ݗ@��%u#H[9����EP)�rF;���;=���@m��X�^1Z9Q��j��v�`qc[`�,w���+��Y���	�B���-.Ъ�[-�ՍV��3oos���T��{��Y���誀�l4�T�+tN�����G��1^Œ���sb���eO�`�,��='��P����aAd��,�ց�A��^$��RID��z�,>��Jht9BɋW2Ѷlo�]{��fkd�����Υ#X��6r���Ϥ�Xjn���`4*����\t�l\�όW���8�,�F�/�K�����e�|$�+�坏F�1N�;�"�A����2�"DN)���1i=ѷ�d���1�סZhv{���vǩC},Ze&�Wl1��� �ECA�话K��B�/���p�x�#Tb*��`X:�  �F{=��㝚P������!$����SL��n^�,�up�m#�^�t�iS� B��Š�L��; �9]Un�TQZ����Z��I�=�N%�c���ƽm�}2�o3zo���GY�B��¹��S����v0���Z�Կŕ�  "ױ*f(�c!�o�$��~�|�P�?�������D�u��q���Θ�a_/X�~�4��SAl�%N�S���[h(}-j	������ݯ	$�Z�q�;��8��d���,�L`W�J�$2$���d���?�(T�o��aJ�����jT����Va.��skv��Ĕ�}�L���:�y�P�n���eE��ɋ���}|�=5��P��#̖��.�?�L�R6���Ǭo���Z�JF��ɢ��M�d]���N8�[�nC��*�~�����@�����N.B���/t�gCR� P�!n�,|wX�_Ԇ������P�i?���U��ە_�{�3tٗ�=�VEի�����ZW#!>Q{X�L�7.q'�F��]��8A4��ow��3��g8K����W���~�ɥ~�
 M�8��k���թO�h6Ti3H�%����#|<�"��WI#��͙8���-�#��q����M2�1�e�*��?�X�g���P=}�x3f���H�:�βu�n��?V!p������hB��ߦ\ϟ���F�;��r�T]����!b�R��a������I�t�����+��JN�oP�w���7�@D��(�����{/�j��{�o9\�nqe��.O�9�獟
��Y�5�|�®����M�~����|,Ҭ!��h4��қ�g�F�rȱ
�U�W�T�P���Q��J����,���.���|�{|a5Vx��v� ���<�!�h0�eZ!&���&=Ӡ����y��
J'&�^YЇ����b�f�(AR�jq�A̘ǫ��,����
�:� &hk�mA�pa<�Q3G9V�0Q������V~a2�$(�fue��ȸ���{e���U�+�M�f�A�mO,�W��f��Yy&�$OT��A]�� ~{a����6���#��7H^�ty"s��3��L�,� BTɈ:�����B�L�l������ʰ$8JUFnD<<8����|�X�]S�E�keV��8h{1�I�N���?����jz�W��Ճ�1ᄣ���pC6D�.�Y�h^��PՋ��N��IuQ�(�c�Q��ݡޏԹS�/-�c����H�NF��f�Mha �C��kP2I��%�c���~g�Յ��mx;.�{uA��0��O�d��n����-���@O��Y�����㜶�
�ܼW���'��&t�;��j BгF�*�BtN'k��0+�\���^�"_y_�a�D$�?��+냄B)���e������sq�67���`�]���]\�`9" p���w�$��<�P�߲z��������쌞�7vK)��q(нN�v;\}W�|hsL�5��9Sr�dw���s+jx(���\�JgD6��ބ-����Ħ���״}��oz�r ��8yɛ��b?�rf� W��n���w��'jê��>MH�{�-�9��r>��q��
'\��W�`�-��=?�G�4�Z� `�����4�|�$� ��92ܧg�hB&i�e<�Մ�6rF�q	�A�셑�0i�-m��?��V�x[��Y�;��t��[(�\-�d����d*��$�,��y������T���eF'��h���;���1kI�߈jS�"S=�MK�T�&� {�&9��yI4����ti����h'�ftl�.��q�f���Ü��IS6b��~UP0�@l$H���i�V7c$�Z����K���&������\! ��ٔ-^�MND��n�
G���wQ)F�%�B�A;�I����A���::�[���0�"��ô�S3J��� ��НLb�[y@\��:�*R�gzxE�'�kP��J�)zl7[�l@�	��x�//hY���4N#���,u�/J�|�5��v�Z����jl!p陖P�����NZJo�س��cT������7,�;����~z֬��t���ڣ��FV �+{��Tp�Py��?Y�5&H��D�a���r'����^����G̑e�� XZ[�Gه��ak5ԃ��di�/���t��k�	L3�k 	��`���p7�
��뚙��oJ���h�>��R���A;]�Q�K�I���3R�
pz�}���kB1��3�CE|0^X���:��?b���@�wl�iM ?V��(�f��M�3��;���� ��ו�(���ݒ�*�y�+jfj���ɍ9⠱��䛔���{6L-���I=Ba2	���E��ė� \�yh'���� yU�Z_�t��7w �\'o�4LXs�i����u5M��6[V�� ��m�W�`%��SM��R�;���v8k��z�s�1R �e8֢ۃ�3����	z�.i�c�y�>$��V��!k}B�`��e�3�5Y%���3j�U�y�Kj�W��:�O �"���7j ��-��%�b�s��i�̴�愗M���y�YH[=�rv�yxV3m�����F:n��`��x+u����u���ɼO��%c����-v,.���g!�	B��L��

�~�z¥�; �^�d	���h>*�\�W�����l�QU�������W͢uN��^�:Hvd�*0������C:Ea?�(SY|%�`�J�質b��g9{c5�EkQ��Xq&/W�,�����a���D�i�ۑ>C��o�I�(��O=TV��W�����"x��+����������LϜ���ef�v��=����>��� �x���q	�B�v��ȨZ#S��H�+v�=Rg���\`�p2�f�������kHD�Ӓ흞_�47��FZ�v�2����V�NS����u�E_�*���R�����"�`�Pe�E��� ���Ҧŭ��)���o(P���v�5)��SD~V�eU�Zb2ov�3>;i�^w�Iƻl�/��{��L_|�Ϸs!��VEP#qt�f�����k|�{�h�����va\Jhs�`�������0�l�ڢY?�7)�x� L���R���J�-�#���8�A�1�
�g�E��~�u4~}�dH�>[�[~"�E؊����>�n�**�n�P/P�4�/��^ys�O�j�ΡA7'�Al�-j
�Q�3�6�m��dԎ��;�]�|�ǈ�^���h+�n^l��tB�}�ݵe~`��|W��2���
c+���G�C����e���i��C2�$��v�@�|�2���v4����!d�Պ�<�\c5id�Dpr�]�'���\s��j����Ls����h���$W�{�)(�2��ۛ~������6fH=Z����D+U*��X��gu\�Z��?eq2m/�\�	'��C,qd F���m������Z=q���'D��S�x�]��6�b�-A�̰`[X��p�_)�S���C���[�_�rOJu;��Îi��;��hH�õ������\���V���]�:p�;IktXds��ep�R�UZѩ��������D���L�k���Dl�W�g	���2�n [f{XSgG8z]�Mm4�+�Fh~���ǐd��*��V��^Y[�@f=j�hp=h6�'6�|I���� T�Ԅ�~�#p�bBa�{�hT�n�svo��]�hG�#V:��v�'��85˫y�6	��K6�*��T�G�*��$���o��Fa�:�ح�3��5��kc,�s�3W�eH�Z��š>N��@�IX�����e�MWA��5C{�l��^+jNx>�>[@PJ���j�]���vީ^<�G|s�%=+�»�r����g�K�9��,ű-�U)�6[�R�����������p���
��ʇ��iq/�#��
�[z�&_R5�w-���{����*�&̼5@~�zގJ��	7��ޙ�hi���nP4�=��S	�J��w�-����w�w�Ĝ^8�&b�ލ�D��ޔ�-u�G(�L��>Uie2��r��<�֤!�Jm�|N�]�΢NC�q��o�*��Ȱ�!�9���Lt�[����B���ua�q9՟�F�٤�B*받�-���W��e�id�K:��N���%��)��֪����dk'U��D��`=e�Fr��1R�����vT�-�|��R$e��Y+ ���4��������$����m��e�?�A�x��ͳ>D�{�V�w�@������3(��� !�N�w�p3�v�0gi����p�4xa���b����аu��F��Z��J>�0�FR0p�W�!�����BE�u���{+��0Q���f~�Vw��;�:�f�]����*P���P��_\�X�,x33G[BɆ�`ت�$<�켷l�3�_��|�L������ �G���Q?A����E�Fq�"ol������Q��Cf#��Gy�Z[�����# {V�i	Z^l�`���T���L'�j!�e�����_	UP������c���t&Z�w#f�@`���y��n�������"M2x2��Z����ۃ��<�%�t��BA�����Y察ɶ�5��JH��=� ����
 �3��m�p�-^w���s8����Gʎ�k�d��(���۾�m7��$��O��Ĭ[w�^��C���� ��7BP�_���W*Bғ�i��G�h���Xٰ� O�����%�U���.}Ba���\��LE'q�� "��,~.�5�g�N�o�*V�9?��h;"bÓ1���ϔ73�d\lQ����{��PD�v'���۔��2o��f��
u*�N����I�B��������W��`�=>��2�p��r��!���s�o��������_K�i�Ϯ:��K5'Գ���`ڕ�q @{oA�X:����M��TL.^�9�E^��\rPI�>�ڶ^� ��4�/�}����T#�v_�@E��o�N�X�����}�,���XH-���?����k�v0f��Y�����}��X��?�5֭����X��Y䩊��U��pdwކ_Q]��dl2j�67<��Q�;sx{x�|ȌQN2�<�>:�D$��^5l:+����c�Ý�}6y����V���q�>:�e��*r�Mn��$Zc���.�Epv�#�R�5e�����3�o��U��ez_�ɀS�=��-��qOD���?�w^�rw�ƺ��kmw��Ht�ƈ� �ͼ��B�b��1�q��B5{�@��9���a�E�y.Hӵ醞&sM6I(�R��D�:�����vJ�wo_2�Ш��nz�,��j4q
���c;bm�'�����1���I���I����I�3o��0���Jɭ�򂲤����7�I*C$�������"�Y��csg����>�1���lW/;���S6���� �l���#KP�ŗ��#�ڨ{ �Xo�2��|2
�����:-[-�2%D��z�K�f�2����|��V�d�O�,��(�|�`l�fkѧ�K�?�d�������:�>����i� �j�A�&��Q�TV[��|Da'C�
P�FR�'>]�
��Zj�0C��2�׎�kX�J��C�v��#N�لQ�|_n�DL�}�.�#��u}>�@���_YQ1�<�vڬJ<���{���hV,���g"	��>o��)�";lw�|"1���üt�ȭU�S�yB��[��5��;+q��X�t�����n7������%U,sp\������x[�mC,���\�W��~m\����M�@���8x}�~oi����6Gs��l��fG�L�xIQ����X�w�Ho�ز{f�<;zt�
rJ<1�f<jШ�onl�F����l�
��D���e�j�/A(��tq<�Z
�����qqC�*;`��)_!\_���_}��8�����C�>d���U���QS��MP'B�s��uPjż�q��:�d�7;�[v������M�u��a�����ŀ�^=�U?Z[����
[���Q���մ?sggiͿcM��)����)��]���ˋ@j��B�4j\��v;�1���Tí	I��Z~q�R����'�̍yj����?/R�� ��+�=����4��U����(D>�J��n���T�k��}� y��hcföJS��O�t���X@/q]��Pp*��.(�`�ɢ�X��٪�b��iy���H�lȪ\�&��\�c�[�C��Y��M��a�P�U��1�-�Y�c5���p?�T���e�Mɉ�~�s,\��(70�W���<��>�V*˥DR,�,)�F�sP=MTٔ����̂���#����h���]��ˆ��Y�J7�甎��)�)�<l�� ���@�Џ7q?��5Eo��B�rP*H�P��B���:7������NC����8>�y�]�J�#�ޕ{�%!_�W['f�8��M�-Y�j ��㶴4���*�����T��|�^�T�s�3}��Iݩx�� �/�[d*[�BT|E�IL�Fb��l��>����,t��C���<瓠Q$E-������-z��=-�e���*�c�2�Ph	:9g��4L�fw��&U���(��4�!�0ˣ�O�Z��j���O�DG�5���4l�n
��'��X���s����fa�{������q�V�4!��kP*�����?�w@b�s$�>����fX�+2+��[Iq���b|�T�� (���Mw�8��G�=wŤq�s��,�F�cK�p���<�ݥt�t���˷��Ƀ��I`���T�h��a����j�/l��r�ԇr<���حvRP�ˣb
�v�7�׮1؞b�CGz
�W�4��v؝X��P����.IZ��3_<j����xt�e�����j�W@T�~̚;�V�J���f;"�Q	>��h��ۀ8�W1��� M���q�|�8��>��FX)���& D���9���l���%�O�����v�F�Or�zǑG(��B��ո~���H�Mko��W^F7�{�Et�85W �uq��ڀ0ٲ���*۬s�]*<&<�~0\`�j��x�ٲ��?�Sh�-V�,{�w�P�wh�A�ed���i��?��}�G����/�Ύ,��O.ػ@�Զ��,gō��ٜ�kP����;��0�"�9��RL껷6w`u�����<�v0�ƒ�b5�q���@'[@���GV����_F���0���\�T��q�y�d؇� ��ۺ����l�
*��P�|O�c��&Jǂ�|�=���&��Bj�x����x��Z�~�"�v��oy,\F9hq��@z�f�h��l�Z�H�a}��&F1t� *(n2��R�Y�/�ȅy�t� ,,=�# �к@
�=U�f��j�bǍz X�Q@��T�FR	�Ji
I%$)�by�1x�\Q�C30�e3�y� �wTŅ8z�m����:�j�-��?'�10�eex�{*���	 c�������c��7���Z��uv�Ϯ�:>B�����G���]��0L]@;%r�w�!q8�V��{�s6�t� ���!��ʦ�T�
}��vR�L�;O���>n���j����~�g����>��#(��p��1�4~�5"R���4� ��Ǭ'���nhwď��D�+W#1�S�VB�z���s'��������J����	�����i�BY��Ġ�i���n��]��x���gMa��e1{�P��f�ɓ���c�i�7����"��͡ZƢ5���ˈލH�n��A>_z���0N=5u8z���P�~�L
�������W��(�{�a-IG�b�S�!����0auNT�O�z��j����pNҾЉr�u*:b�o��gIѓ�e��,�����Y���`D�9�:\qS���ղ1wro�gw�t���C<ic��cd7�9&�D�����RUj�f5o���< {'>R\S�)���w����;�"T^-��w"8H��D2�)�I*�{J]��	�n�efy��{�oFL����PW�kN�-��oڵ�9��lGL�א�5G��+��b>�7&J�=Z�NC` ��&f�_U�<p��΂cMTM��� %����>�M�B)�&��RE)����0h��>~�d1`��k����񑂨���r��;��Q�_~�&;==%敆���\�w�QX�������f��l5�U3�Z��䲷�N��:�	�̚aRb<aCI�.y�[>�.�#m��a3�;X�W$�Gܩol�-�L9�i�Nc���ql�*�Y:��?sI~�6���^�פ=�%���Q�A����E�r��k�U}9YL���"��^��]���:��I!k���~|z�Xq�x�&��L>��z�S;JZ�q���x�����?�bf��K6�HW�D�|�ޱ��D[&9m�Y&c�r��n�H��������m�� �|)6�aX��>'�4o*Ћ�����6Yx��)�a��k��^+�H�[fJ���uQ]`��a�� �=/"�p~�M��~����g�4 �Ǩ(h�:7lX��L�ː-�pP-�4�h�d�I'�>�ze�wo>������������ ��1���� +!�y��lM����̮����0�8&Ω��*��<��Dާ�ZN�� {皹�`���.��E�O�lY����c1��a&�\��1�os��@fo�Or��x�z�S��� �K\R���S��l��X�L/B��x�[��p�1�MvN)*s/m�7.=�;+���Nў��m�è�m��6�YdO2A��r z����%[�AwB��*���HJb��G�;Y����Yj�m���I�Ÿ��g"|�%��5D8�J	��(�]�X�-�&Q�1�騂��e�㘅Lc�Ա2&�҃��?�[|t1��~���q�ȥ��SY�7�ܩΦV\��8*�bv8c��|�������7����	�J?�x�e&�	9���A&#��&��k0�;��i�Dmt-��L��nO�b��"���j�"�1a7\�D����E�C��Wh�E��_�7j� 7��=zF|�}���$M�c���e
	�s�����J��B�k�J�gr��E@���O�lmw.i.7��|����K��`��G�..��l�r��z$�Zl��<��A��M�Ćժ�h�9�)�˱��!yΖ;�����ǲ=`4�[C�ҚuPuX��E7,\�F�t/���we��r�7.B�2�ĸ��9�%z��x���pmK-X�@	֌)�]R�!\�yj�4b�*�?tH&@S�{o�VCG.��%��f5�J���`iC��TY�_��)�Bɿ?���X��$IR;��WnA�%��緉S��EiTl\�=P|\S�\K�����yՁ]`�|t���`��I�P��.�=�k���i��"(S�s5
��9^�+﷕*�N�x<.5�o3�?�#�sgh��U��,p�J���=�)�6�7������D4>�����J%��f@晜�i��3c j&ZB^�(8Eʢ��a���-h�q|-���ga�d%�s��jRvV[��b���G7� ǽ����3�1�����j\+��Kn%G�x���c��F�}r�\Z�+�~��
��U�G�]���k��� ǅ�~#�Z�����D;�c�_���I����-=���!{%�B���C��.�r+��(�����A����t����H&��%�ZQ�KH��ڨ, ��y���WS�!UZ���6��GX�Bs��Y�Ij!a��_��g,4踝,�(�r��� ��fD��2߶��CQ���vTC�M�oo(��p��_ x��`����F>�s}��<�ձP�^-��m�򝽌�`���{^����Y�{-T��\2��GH��v{�y�n���D��_=��]� ��K��'Ͷ�p��7j�OF(>A�>���uB�Md�L�w�3��I#�F�Nēa�+�B_�{�:N�o+b��֝��b��,��7m�B��n�rA��`2���C����F	��<����-�Q�����-x�!�P�QJp	����TE���lw�g�=��Y�ߦ��e����3J�u�'vEJ�pHFm�l�°�)���&��̛�h9nY�"8��ߒ�T-L��U� ]I��Ȼ�m���Q2��\���S��C�������&���H�(� ��˥�� 2U�@z5�V�!��R6jD�v�(���J"��������2��Q��l4y��g�����%o�W#P����4-9|ⶅuw�J�hF�W���L9�o)���R����y��"ĳ�5�؍�П׎0���iЅ���6s�;�ӈZh4Bjh�M��Щ ��\�P�2����.AP�\�u�e�d�$HJays�t΅t�H��Ǡ.F.���M(�ޗ��1Y�lC^AH�8;/@�]ߜ����bi�S���µ�#�/ʴ����l�K�qeO�5G�����H�F!�)�#�˺�tPY.�U��Y�z�C��I�J�F����� ��|�Q�1���k���H^4G�Lp0�F���.A���g��w�
C-'q��/��T�%����/��D���k{��f�jC%G�P]�cEf���1a�{�0{}���!��"��-l��6(A��]ezA�����gAT�p�x��<��N��kQ��褡C��g�K2\ސU�=������5�V�HJe��E�u�B�|��ф�bN*�L��5�"kO_bC���ˌsxR�ַ��vV�D����Z"���d2-�:��Z���.&�m���7w���(���LE^5���5۷�۶3�׽�</+��HZI;��!B>s<oH�.d���6� �wtQ�<�8�x�Th$6�9�ez\&���q�).�z�u/���Z�F��hlî��.�o;�����[���@�#�/�z�p���y�&1L���;i�{J��sԿ8�D��-�˔ï���M"�8������h�_@��z-!���y��H�#b�?�rK+;{��ƍr�=�7��:$��}[g��SӍ����u������A!�a�tCu
�#ɀ��Z4����HG���_�Yp��Ɖ\̗���+�X'������ⅳ{>��Cyq1��md1ѭ�>�O�E�_y|X"����!v5	����LuI�[�[:HAs�c*ۜ��~�M��ˇKR�<�S,�jSA�Yj{.�� �Wd���X�&��e5���.|,\�hTD;�(�c$��?�Y�(�H���iWlt�;aZ�I
�r$zp�/���'��hBl>��C��$P�2S�8��x�M	O�01�/�;��vP���4n�4�%�(�^}>��YQ�l��{��HA������Rea]ӲS��_)Q��k�-b�$K] ��R����?��N&��`X�sr�h̃�����X�$5"^�g����Ʌ�?y_ذ�Kꐵs[��/xqK?�1��G}
4t����Ą'w��K}L�q�E�H����T{F'/])�\5�1��A{�F5/�e�V�
.�G=��2AXP����ĀSK�G8_`,��>�v28���=4��1w��f��& �� :1Hc��	o�������c�O��gӨ�@��Ẁ_�PZ�E)��P�T8�lH��G4g3�j�|�*� /^ލ�;ގJ.��0y������ſ�3���9Ӛ<�C.� ��?[]�в�
��=*N`?`cw۶DҕJ�
M�����6�K���*LX��N�Ւ�M�,!��T)e�1 }@�d)��Ȝj�ts��}�0|ބ�"c�iA��k�p}�����Cz���D�mU
���ӁO	�h�����i��g�i*��`�l�e�vݭ��[~r���b������O߹�>ht���TdD���#~���bD
�-\N���x�u�|��ݤ" d�W��Nf�x�������y��'�9;��ȥN�n����-���PV��cV7ݴ���@��ǙB��q|��orR1��~���0�I�7K�\��uo1g��(Os�~:Fp�A����^Sp�x�e[����L����^k�6��K`��1oc3�c.�(�-2G�V�(��0��-�C�R}Dԡ:FI��N����q;�=3Ŭ���D6kB_\����n*��G؂38��W�]�xJ���'갏����W�����Z�uD'��Fg$��h>Nv�夵O}������et%�ʱ��<�Z�T�&K�8�)��S������j��Utm����WNd�mR��V�<6�z���ʸ��K�V',@� ;� �n���C)1F��O�s�ѵ&�H�,j���rU黮�Q���ء\�Yy�U�;����J;���$�pQ�p����@H��٫A�BՊ����rjd�
}�9��t)�0�:b����?�vJv/T�"���k)�#hI��\��L�Sc]'>�75;�E���c�b
�%����kS?S&�N�Y�C�
&�k�ov�R�ʲ�CL>-�����O[�r��fFٽ�H�^�ES���,���y�^�]�F1V��5��mA3��6��M�\5;�%䌃}i#b~��w�����I��_���zd9�)g+�*��s�7��(7o�����&*��W!{��[���ֈ�5I��'�5�k�������NR�֧���ȸ��K�����e���q$�w���֮ۢ�WN��f8٫?}��-�LTh�큁/&Z݅j�k�=�����~>\��
wkٯX¥���	���^�=m0���l��v	9�;LO�T>�K��^Xh�`}��^��l�.������k�0dWM�g�O�m-aG�5x�� � �촎�|Q擺g�p�o�͎G��0y#�t�	
)��S��[��(J�(�qX*��f����Yje��mm��5з��k���]p ��rQ�.rM<�8"Rx�ia���%(XMl'r_��W�e�8�m�e-��3!M�[ன�j� �ڸs�4I��k�ў�c�<c���i��I�����P䦤/*�=�4�������o-K��B4""e2�^��u��鱯�J����g5�l��4��38n:e�Ⱥ_��\x��5�ҷQul�qAgs��I��
g�\��gA=
H5�� ;[�e`Y�\G>�xP1�Qz��9n��&r���L��zyo�B���\�T��j*'3,�B��}���@{L�����'�ѽP�����9#y�ۄL�D<�]N��I[%����YXE (��������'����ʚ�2Q�B�A���iʠ�M�![?����3~�kg���ZiX�;�� �W��8]���?2F�u��
uy�Ŏ�K2Y�Do��x�Jm7�{0�A(�ۙ[%��� 7.�����ˋ��v�ŕ ����X�Fg��U�JT�Xdx�؇��7@�'�Sx��u�RU�U�����.*C�N�򟠍
�����#��ɚ�ܴ�Ο��'�2j; ���-E����=�{m�Lm��2T�@���Z��V���뢔}��;�6�T����Аr� Q� �t�X:�Y\ފD��Ȥ˵�{�!	��$����F�����[���X�WI4������w���Uxu���~�@��Ȓp��ש�����*���P��.|[�#+�U0����M�[�4�0�V��o2�p����}IwC�~��Bh��:I�ҝR��.�۪�𖅨�[���<.ۊ��Zl	��*��Sc��4���#�4W�K�u�� X"kC�H1�&��+4@�ϓ��;��b�S��/K���B�����t�_v�:l;���)W�����#>�c��cWP�#�%�aP�{�l��"{���T=n��xT�D<;.��ۚ��#��^�"8*M���p�,�B��>�d�w�	rU��$,DP���F��۸��3�{քgĄR���s�~�w5������i��ز���˹٬^5��׀��t�Kt�|[��)6��s�	��1"3@1^�B׹K|+r�0��t��M�M�gU'\Ċlq 6�%�_��VM��ǋ�&1Cy�axOٹ�b����"S H��=�If�xi����d��PM��0~��`����G�'ͻ�˽Xye�<�m�?hWN��pB'��^(iyc���%�۩�M�Z0�׌����wgkQ>���h�Ѯ9Q_�6&�}���>�3!��b�nFB�����߷���F9p�'��W2���doVT�m����fd��1��V��3`j�'t<����k�a8K-�E:�Xk�GU� J��\Rzy&R�"q�3�0$r��~�̡|��}��i��"^�0�s��fC]�Y�R�!���P��B�!+�
�s��ӭ���n�I��[�rVH'B�{N�%��ȭ.�˭�"ױ)��wo�ɠ
l��CAY�̴���Ȩ��;we��LU�t�Y�c�tƆ��S7�׸��&�ۿV(_D��㿦L�7�ʁU��3�ߚ_u�+4B�uA�Q����x8.#1�u����2t�N�Fv�*HӅr���F�*L����sֱ+g��l�������8�5�]�` 쑙"��$�L>�/B�M8:�%u���H���Yj���C�(�N��בϚ��/��p.����ؒt,��q�h�0�H)Q3W3��|R����*�$-ȃ�ҥ���V��>j���9qlG�U3�>ř��еA�#]�j���3*gEs�R�>Q�3Wٔ�QI�!..����m����<����}���֐6��~�6ڴ*��s)I$r5��gB�Z��3)�Jht3YFk��X��{[er��x���HF+R7�Ьd|�Q%~z��2y`��������ɮn�����7���s�^dN�iw�x)mn:��� ;��;���L
Bo&i=_�����<�JʈO�73\���E#޵�Hfj�5p5���z�LʥH'�W�@��;n{�uQ��4��g�U�$�����罸�����~qǽ�zz�����\@ke@�z�� #�4�;��Y{�On���[��'yB���A <j����2()�|��}���#��~��Ϛ:
,8G���Fu;w�i���A;��^�=
�s��ƶ,&�u�:2�`w�8xh�����ez}�c67����8T]����� ƻ�_�X�y�.�ʥ��;.&��1�6.|_zw�)+x�_Iw������\�����}��L{"(�����ah��&�95��z��Q��J�R�X����M����,{�s�(
0n�@M�5�FT�v5ᖂ�?�i����^f+mE)�.�쌨���6l]�Zk��jKЀ4��1�l6�xs��'KN��X� _���eh)�Α��Xd�D���u~uhl4ZАˬ��v�OM��Þ��B�i�ȉ����!p� <��֟����� ����B�(*�/��	儩Rz9b�$u�'�r��6�3{�,\�!ȗ�/R��J�b�ǅ�"a�ҏ�z��?=��Tܗ�=���9v�@	���!:G�Y�<B��v.T�jpX�v��H�~����� �t�����^�W_<^w%1�o]���c�_$�1�$�I%�I��ha�Kdۦ-�3�
�������߆��5kb����Ӂ��,�9�5)k-m>��x��!��;��p?�/��\7^��!�ɿ�f�u.��S�YĕuYX����ˤ>N<u�~]�Uf7�:b�BI�8����?I�p�!�ϭ����ćt_<VA:�hCM,^�J#k�t^񢔶���c'���*0l8P��^a"1Q�-Nd��fꯔP�e:�O�0	��M<�'��Z��L���&o�8��fU�����(���&-�*A�X��>�ÙPbq���}�E�Hf:��~r���UghZ�.��;V������ JK7���8�Kة�8��{Ŋ��tN�0�mL,��\�8�4����C[�2�0=]`x�]vw&}����ShPENbD��7�?�%�ϟKP�Y��`�+�f�!�r��(����_�N�3���f���퀛�÷/8^D�7��Y<dw��|Ȕ6j�&nR��>���ʀ��0PFA,�5$s��:cpd�G;^�kY��K�G'�D�a�v���L�I�SJ�C4��3R�<\RmJ	-�G:���5hHt�[�_9�'~݅��E:m�4�>l%߰wj��ς]3��m�V'a��p�Y�Η�r�D	��@�G�V�F.�4Wh17�=��k������5�Z?�w��2\C�-�c�*�q��It�Wy��I��ĉzW[�3O�"����J�LO�kC�U--��g�!5.�E��@;���V,E�����%0�^{Z��~��������,6�ld��J��_J})Z�C��4]zo�dY�Hz2���~� ��Rq\�-�A�ѻ�m���;)��*��B���qׄdrхȚO��4�]��Ȕ7�+��@�tO�s{�e(�&�tɩA�ΔK��J>�TG�e�D)R>���wP��bC�-'Dڝ������,�z�sͩz��+��Z�]�C�;ˑo��<�A���P�k�8]�WH���/1�6���(2+�5\�N".��kH��GI�������`�cp;3�qh7�*���aSŸ���c���܊���[�w;n���=�Hp?���.�̽]�B)�~����ۣV�������c����1�j5�w�z�:KR"{m���<����#���?/�La�[͝,��|2[i%N'Р؛�RQI�+*�_�[*�R=�%��N��" �I ^׈y��<]< ������E��_�r`]F��So�|�2	��Җq8n��pGD8�T
�1L �jo~����W�b���Ii�'נB�3� ��Xtc��H�9��� a�S5����j��a���ɌFVI��W�ڋ��*g����|O�����Nl'b[��ƫ	D�=[�J:��P�nmM�j(����%��K��sQUn��"�w"���(o��iE��f�*}*�9H�,+)���O�.��� 0�!�(��Zʯro.h@.�X9c���w�$���\X�GӆK��%t�N�^)^��vi�(�=n�,�Q�e�E�����gs}"���D�џ<����?:$�����q&+��|����K��vr���EZ��$�buưBÎt9��&�����J�]а�"Ya<a�=e�#\%LK/������b�-�hS�x9Y�+U?@�'��ؼ3G�$/�]��>�Et�S��z^�'Q�C��?�#�&�U�2� G�X�vY���zò᫶�s�ƿq!9��5v��-��vo�sa#�!϶G�#��/�pB�k c�
}�=�|�iG2���Z��8����a�R����J ��5���܋d����.�B��P �]O'*n��c�� ex�+☮V�^�"��l\[EmF��G�}-�(��T�E��"Q��b�.�RT��(B�/1#R�<��B��r�$�:XKf���=[�N6�������s�Ҕ�!��EWо.O���!���Q��ZHa�j%�t�\*a�y.�귃3�7-�PY�T���D����G�B���\�w�ޤ����F�3%��f���瀨�z�	%~f�Cf|�C�Pv,�W{�}E�1�1�/�͑U	����5���d����t��8Dg����d��0�hY!&�kR
�c:�*�����o�{�j����.^��<�5��>x��u��F�&��[�K��o�׃1��?�6]ϩUI����'o�y�=�D4@8c\8����Q!fm�T`\*]�`�U�@6���zN�mf���������c� ��a<_oPp��H�Wyqe�^9���)�C��S������\fH�˲�@2V��g5�!]��Z�=��,r�O��^�ݷz��40��r�=��Xw�}�����jyn�f�
jY��Z���ĉ��a⻜X�R��Z
6f@�����.���}�{����]���5�,,��k�U �V��t�5����Q������^K�N3z�B��J�j�8�}��/�<TŊ�=�7k$�~̂=�uzV��ϯ��om�����:lRX�0���>g��wc���+T���� xY��PF�9�I��j���m�G��6�Y)G�^�74��22��R�~�q&N�	�1��I�z���m<��(_߻�ZD&�I'��:��?u�q@�M�8zs�Y��Qi�F�9�͉9���|��[��{�1+�cY�$�w�hD�`x�9�o{7����=����G4�{F��L���@XI����]�ʔ��������U|��M��%w�4��*��f6/���N��D ���.�E�Y.�ѕ������͊eHy���3��e��¤��$ N�����8�Vپ�5��2���,{���E�P��"T�*��1`LJd7�t�C���B��>�Ԍ�&������ꚍ�J�+n����Bd(x��Rk��λ��6�kRo�i�l�5R�N+��&�}�2Kȡ�l?E_��d��*P��h��؟�C��7�z��ThxE�Ŝu�S�o^����fL�U�@XY��2�*�œ#�O)	��ǁD��gf69]Ы�"�!z]���K�k#�)ZE���k2Y�7A�z��m�ӹ����gs�5������ ]�'\�`aDsj<�����1�4a=
uʊ�3���F��rdt�����j-�s��mvQ�fKs\)����h"�\?���g~��f��z��,���A������?ó>�A喝]ࣱg~��Lv=*?s� #�ˣ�i���#�?��)|���f��)�^@��ͦv2ܚn,�k��W�#ӱ��N�ވ_�=5/0= J��z�}�o3yK"W,����7qzQ��!�2�+�_�8I��n���?�\�8��
�뮨���EԤb.�L�%��+A(�g�7a��P���X�1��27&b����	հ��`� y58��+��$`�������s�O���୆ -�}�V��.@i5��[z��������Mp67$I�vY����ǯ7�5�58��*� 3����")��	�-iTyѥB��v��nG��&�β�7��ϣٜ_,+agM!]:�`՛j#Hߐ�O�΄y���=��i`-I�Hݬz��@��])㪶f�6�PNra�q�,��.�}��إ������'Xݚ���w���m�e�%�W���~v8��c��@Y�� �J�%��8�(f�Xi���^kĈ �*����I�d]|H�G>��"\H���T@�b.�}=`C���/�20�vt����s�]���ۺbL���_pbҋ����g5�#GF[�c�y������)���/	U��S�(V�Q�� 6�Z�lc����R�x?x���Z���Y��B%?��i���ad*��-�\��8?g-���'L�FS�\�d����=��a|�����N�E�E�޵�I)����=��]��^��+�FO<�?J�aN���
Έ
�U�V����̎�+�d6[$keJZ�nm�sZ=+����f'��w�>w�a�a���'�n��/m�C;����Ȥ��˵�V���K/MW�%Sg~�4�~�Hm�o��r�׏S���@����oS��H1������ �Q�u�~H��2b=��}Z ��K��럤٬x�z��Kh�͢��{��	E��=I�n��L�tT�6��"'7��j�!)���m�'��� �������l���#Y��b�u�����w�D�{���GyHB������+��z ��Tl�#`=mZ�O�jMؚ`0���eyq[��F�R��N�旍��xYQ9$"�ڹ3P���>Z#���5�wWj��6K!�$$)j�&�.� oC7��|�����)2�%~��"ra��� #0~����6��]H��2�	O�� 0�9��Ϗo��i��ߋr�(�4���A�q���p�xN��.�|m{.n	�X�Kؽ.K��^2TL���刳w���1���(3H[7�	��+*���Y��s��-6�L�f��<�;O����=;5��˄�r�B佒vο 36��C��qL���9)��*�,z�O�T��X��O�4ӝ;��_�-����>#��S��Z|������5ئI!��Z�x�aF��>(*RU����cjiX��
F�@��(iؽ�rq�9�\��F7D���8w��<\*��;R0.��[ �s{��R2-@A�1��N'O .;�[���Ihv!L}u$gp*���O��:�p���-��6���.�G�E��V/{�Yi�i%�/]ͼ��?p�v4�I7���
���0�c~��&��r�>V5�v'Fu�y�5_$����Ñ
X_�l�WA�3�
*�Ox�Q�o��T����4cl	���MGS�Hv�F�`������%W����kJ��R��զy�U�$>
5��z�߻�e�y":CLx���W��R�����gډb���@!�:�E6�S���)TQ}�D��}U`ɐ�t_���#m��������)%\LuM�+	�t�F�;_��m�x�1�P�,�!��^��:I� ~_`��v��M�Q�?�T	p��U?yE���p"��Tj���㱇��%VƼ��L�Q������{����XJ?�������{�0o�I��jX�u<�7l����z���"4�ǊA��_di�n@h�v��1��7Ք�����b�{����v	���v^m���9e���e7��ȱ���\�(m�b8A���L}���̏J��H��Sp���s��k>2	�h�N$*�7�I	�6�3���
�X
�i�`S�X����ϩp��d�Bt�o��j�(Z�Zc��Vr1=Nr�Wx�즌����[�M�d@v�&~r_���u�gV���yIF�q�1C,�����5n��Wx�5��M�Aܕ��@}1�#G�D>�g�ŏJPՠ�5��Z�\WC8[�y�mi��̰ѪG���=��\��eB�����h�9�B����)'_5$6�l~wG,jC_�K���a'�4�sO'���׽�mo���C�=-R���j�L���2��+���{�WO\�҂J�������f�+�[E�^�[��ă�\#w����r��ړ<t
}�#=Ӧ9v<��$���%��<��L׭>�}���ʈ�c�H�~���}��ܱ$m���*�
� �2Т7��+�>I��.Xe�d5����˟	(R�Ĝ=$ҿ�]����;Ut�U�I��+�Რ|�6O��!Sh��.�v� �k-�Lr	��?x�8��I��D�y#3}�ԑ�t�ۣy*��e�<����>���~i!?,b$"r8�(��ޞGK�IY%G�-u�2��N"����լS����`�Zψ���n��H����D-�-0�>Ez�-q::���oNw����M�T�����f�蝲�o��c��#yĂ�@��<�.���r��c"r�:,��w�D�α�9�X6��S{�db,�;Q�`�J��d?��y�w�e.���L����W�:�Wv��t�:�fܯS�Jё�,X7)΀���ᦫ��T�':�T����0߃[�FR9�n+v�ܕ���@kz�&Hu�$��Q	"�(ͬ�9�c*M��1�n<!�&r�6��Wqlg�;S"�wÁ�LNL�������{(1L����Qb"�.!�f�1�Zm*o@i�
�Gb�Sە7 ��(e�����K�^��?7�=�s�6�	d��g T�͈^Y�C��]�k�O��n��c��F.*� ���>i�[��������W3:���*��A^�,k��Q��f���}ħ����]6x������K�γ/D1�Q�ÈY�:����i�͍��bt1a�<�����	m� 	�`�	\�,c>:�X������P���jc���}e�	�������=x��u���o���jV.B$��sG��N7�AI���٭P\s=g�!�wɑZ�M����!����+���l�op:��/�秨�3 YB���9�z��zek78�$�ꦴ�$P�0�_�׮�I̯y3�Ь���"6�ʶ������RTYP,��Z]�:?��iac��Z&ʯ��m��-Ȼ�>�Κz����.���R����v�/�Dp	|Bк�x���Yg��&$�&n���@:��->!8l*i�HD>�b�PM��o����Q��*-��=H���Fn�,>�Y�G�f���4Te'o:��$0�7��;⼯�\ɗ7�����(�<��n�}0��e:�w��^.Ϋq>ӟd��W>�D�
��G捊�#���ٕs��� ����x�CsU�!�w��u��h�T厑TK�A�b.�wC���NҎ��*IG���Α����L�<��&*Pq�{�a�(�I����_kZe�V���"i�I�ϖ/7����<+뜊r{�31,�N�e�b6�r/���J��o8�/Z���r����o貵+�8Ď��'͂|
�ų���^��w�%R�Z�o=w��&͎��M����+��p��FKGIm�]�M��X�-X��b�E�J6�[%ۓ�:�r�Ğ x(�	�m*��-2�ϧ�>�??IBs�jՆ�i�� �8Vv�}Q����t�����`��\���@���;�>ʦ�����s��rf-ԨoZUiV{�H��GF�Ay�=�&d�Y�?=�*��R��� *�b���2��k	��*�v�j�#�_�a>��#vf�'�<:����K�ڣ_��]�v��%ڎ�y��$c���}�K���ۀ�ݙ}�G^�݅��ʀ�_`�3mE2�\b@9�pز2�U�ې���>ZL��=tj9K�fCݖ��SR��u�?]�������?���v_�s���=��\�� ���y�b;�"s��u����}�-X~�T��6�3�Zt���w`=�M)K�&�|;�vC���k�&2^Z�`=0/�~����o��\��BI0DX����}7�	��T?Cg�pKI���Wp���R 	e_l0��/3Z�e�!���/�Z7�{��MX�$�)�;\z<��({H����m�X�-6%ШS��4�s�R8T�����7̀?]O^p�/�[Ջ8��%�i'S��QP�\�2�/g[��F�ƈG7�.�)�8�{C��#M���Ŧ䈡��F����{?ͮ*�FO���K˒��I��K��X	I��:���jH���F[l�ъ�?�d��"�ш`}FL��-��˜�W���g�˪���A1!��G�\��U��R�s4?�d��e=QbQy	NJBV�w�l@{�b.�b`�k
�X�z��y�t�Ӡ��['�t���3�pxlI,B30���C���+����x����������kv���� �|/0`��?x����&��[.���[*��{cϱ��u�Q�˷�M��4����tjR _�!�׉�U"���e����L�Q�6p���O*M�+W&B�܉�dh'1L�2�Y�\+i�mu�c�ʭ�O�dp0LE�.`E�D��nQ�:N}~¬� P
ƎMv{��y	�rw$wq��$A�
�DeG\��x��z�9��^s��dy�!D ��������)]�j9����L��ЂVx>��.�n֪Yu�+��3���嶕�p!B�l�u��I�w�<�íxƆ(���$� ��*���u�T���ڰ�?�,�������
����1���S�BlfQ�[��L�7��Q���T��k���-M�j9mO�L� �kօ���G���k���r
W'��F�i��%��)_t���ld7�A2oА���0�����[W�;/���A�?�O+P�cP㝄��r�YC."jÞ�o"�΁�&�HCgC�5���)GT0f���?��S�}��]�E0�NJY;�����Kl�I�ԥ��v��تUphA����x���E�K�㙅����b���5��������<�s{ *�4cF1#`���^I�e�j��"��;	\t����L%P��M���u^� ��k���gI1\���j$*��|(ϝE��i�A`́�-�@��A^ڧT�Ѝߤ��q�����m�m�b*(��׷�1�����X��=�����@v�}}eN�s��Ë�z�9��;��J�Q9Y�3:�Y��*b*ޯ�y&-���J`�x�w�a�b��{���b��=��C��
m:��X����-�p'��1o��T�g���t�b-�'���CK�B�Q*���޾��Ԫ��Q2d�z *�n�Z�AO@�
y<��x��R�Q���(�x fkK%��ӣ90�_('�J���ą�CB�oQ$�h�0뒑�`u@�lJ��G�N��و��	i�x8t�#^!�!@�CKl��n�����'��N���s�Y�El��
g�H���cǺ�p�uJ�+��^i�"V#�
����X<��ׇ/���ЕC���\��$A������P�Y��%ܤ��;(�cV_ژq]���[Ck�s7sk�z�j��jt��ѱ�d�9�����'*��'t��魿LvqީPa��6�m:���`4���"���	�]@[xË�J�ߝF9@#1Uw��>�� ��WB崴&$����B|�;,��P&Tuu�,�_�%��3g�,��-��Ϗ�XP@��.5fw���P�l�7<!']��+��ZhZ�V��J�Ho����Z�:b�_�S �K��S��&�������0:�窞����F��X4`��uw���10��\��80�ؿ7 @Kf�ʽf�G���	�r�I����S�o��2W�N��9h����ݨ�4��H'��t��#��{1��YѤ:[�<��fb�cy�?�}ڿ���ċhyL�MG�m�0z��̒X;��ݨv�=��D���|�!I6>�>�U����l&�ٙj1c�A.��»QX����o��O���	��|_�͍���5���9CGFt����)�+
�+ <���̷3o�+�M�Zs*Q��s���l:Xr��)[��rY��!��%[Z����V�>s�&dߑA���{�N*�����[�k����nxL u\�(df���4�H&�M���h�6�!�c���b�P��82��HO���#1h@���/r�L�<��Z��F�:�Q�����L�hC跳/9a-]�&%