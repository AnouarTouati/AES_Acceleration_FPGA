��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�
TB�(+�
mQCJXk�ɒ��Nx�m|&�X����!��K���u���?x�K�h v�ag���Dz��ZZ+#�	TQ,��4�*��nu6G}Љ
�2Lw{���.4��h�k���5u�:g�X9���k(�&w�;�V3[ǽ�X\=�E�a��_�K��
TJ���B���|�˥�f��=�kR��ҩ�$�x��v��6���s}u~/~Uº6��&9ޏ١=\�c�}�b<�|-'��F��2.ݔ���l�դ�	2�*gؽ)��n��m�Irz�R��Q>ʜ�7��L����.�n�d��@0�`��'�Oc)�y�(�Ě��ϊ]Q������wŀ�8�%�����,j빌�ت_CeBA��}砋�_���XgZ��)���z�Ro{o2�N��+UV���)��d��2剥����'ᯯ�_��g�x�7�Ͽ�P~�� �uI~�l��0�����{�e��v�Cia���!�}�C���Gd6�����;�/a��:�U*���\ME��pӲk$e�)���z",J7����qv �Z7����=�Q��C���>��b�f����ύ��}���������|������,0;�;�#\��Z)mͶjJ�]�ʆ������Т�m�_�����[���g��
���=]��W��a[d��6�LNn�ɔ�l�jX;u=����o�^vl�����Y���B�O#�Dtz�e={�
;"}iqR�R��b�����p
���'���h�����Z��\�c�,�Oճ��1�lE�NACO�>[q���k�#�{�E�Fre]�����1�L��K��d1�+�9���l�aP��l����1&ۆ�Q�>n���Ͷ��{	��
�G��g�W{��:�ÆYj,3�;pgҪ��(
�C����>$ UDY�ͳ-8P^����sygk�GV����:Y�7Mi�Z�]�0��.y��Uפ�^
�;̹}�1`s���?s�ӵ6��8Jh�5F�P���s�DX,a�f�aL1�8Z�����r�s��7_Jg���5߬d��pFFv���1��,Cr%*t���UTd�J��W�,*cy���M/�)T;	^;J��Ѓi?��/v�b��L��A0Rs��5&�3�O��?��(YzHiOܿԽ�z<[��R�yi('A�&Ѓ����q�&EdW���GM-�9&��Q��m�J|˅��X27�P (X1��hMꪑ�:)�x`~�J^����pj�mܰ8�����'� ���ݫ�
Υ�����Ww�s��%0��oxV�6�I���m���) �F�*j�Xc�1�}�+�b�]I�8�T���Gջv���4.��E�?���"���$�f�dd|wd�v"����'R�9�s4�B�X�B��F#�W�=!!���R���C^, %)��ec�gGP���?ՏL�� M�Ci��8Y���(<� ՝�=�#Y:�2�|;�v�=��2���DIc�:�
�)����]�qߕ�
�B4�����(�X�<��:��L6yb��o��7