��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P��/�͢��u>��b�]���K�_�cx���A��"�Q��pMl�jh!�GC���&�Buԑ�y��WB���{��|-3w�A�#aS	�Ƨ���9���1�-��H1��Z|���>����@���)�dw% ���2�J4��ŷ�|�,�,�L��j�odz��3Q>XCSc�oC�f�t�'��0�I��/[�/���	��l�woy���h�2�
�du��\Cx�io�"6�r%Z�d�}�Ǚl
���m��ļ�ؾfű������X���_�
�	�c_`��\]�x�#�Z�����e[N�1v�b_iu�����m�\%r�K�����s�0�⠫o04��� a$�X`����Ը;�{����M�������OwH�?������;`-�l����2�Wk�b ���((�=��X�~�@����>�u�q�U܅�N�y�p�5���E��L�}r0����� *�8��7������޵s%�G>t��U�j.���7�ou}�A�`ͦ�X�Ļ�
���Ɏ3�\�Z��UF7�+6�awu�ƶ�e��HP�8�ˎ�U��`�sqڠ*���aC��D�k��3�kc�}qҺ|�m* -�߮T�hD�3��s���vL��F!���/����=�d{��I�Ǫ��5�I}܆~�i�W���u�i�Y�_d�D��H�,� �!z��'� �b��Y8]#�M)�A/���ԛ*��g<�̢P�ϡ�Iv�E�:.=OB��~��,��E�F ���q��b	�-�#��|���m��Hx�IB����_C�J��R��6���Z��v7?I9�Q��Y2�#F1���׃!�MW9V %�5�Ȼ�~�'��:�Ho�r�����T/R'
���[ڴ�c�٘7�\�����
�Kp?�'(b�Sw�oEˑh�BB���O�b5]o�Kg?~A�_��2�Z�R�):0S��ؖ�~��-G�Vg�v��p�5Y~�����X��<���R?M��G,�.g�^6�;�f&>�s�+�m��/r�{�f��S��Eۧ��������6Y�����􇬗�5ҕ �X�쵟:VUo~��U���%����F�8��o�Y�����$#��{/�ʟ�K�2�͔pp�]o {��:�)e�w�����=�Q]�{�h��.|Oڍۣ/h�g�%̊�S=ro����F%��;#��T��_�B�0��K��%H��E��*�l�c&
�\��0]Yӱ��ӈ(��s)�L�VEݲ@�ʤ�C�l�:�������()u��LJ��/�������A�<_1W\ ���#+�<�w���<C�:�JF��)cf��Ű���F//e�b�Y�|	˕H��u�����2�
^'گ�:�V
+i���5Y0l����O^�-U��sRk�d% ���U���u��zOntۂ�� �;��	��'TQm�P��}�T�*�K`t٧���y�NqƷg�LV��usb���̚O@� ��5m��������/T%�+VO����ǧ���S� o�+��0LY_���j�Y:���p�9]vш�s�|fh��Jp�bA����W���;�qH8���bg���}l�Q��Qg��wk�0<E�YJ�q�Ic4���W0����r 
�4ۯ��hh������+�b[���E��3�o}#��;fJ�2;J����_�L�N �b��k�i@h�1�N��O�v :(�#-��?k̎<��m��/OyZ�ֹ�}2C����h�8��*A��]`_d�y[�r-&c��?��69�MN�@�l��E=�x*�H4������	�B�=�7�t5�w�4���3���&��U�FlUo�+��ʸ�.Kun�O����<�f��u���?TO܍��	���:m����zwH����R��̺2f����f	c���B��WP�����(sTta~?k����%�V�i�!��Y�U��ƀ�q�d֎R�$�I�s�C)kd8���s࣮��$���5�g�
�M�i�Ә�M�ç���s�)}99֦V�i�B����H�x������.�f����]�Xu��̓��A�;{�� ��]ӰP�,�t�AT&�ߞ�P�e�ϼ;jT�j�F�D���zX/qY� ��G�U"��3]yY"��:��T���!m�%��0܈pi&S�T��-� 3&an�Q��Pe��$=F��x��5��B�ݵVcY�}K���.���r�nQr:&�����o2ق�� �޿���P�T����h��G��7#����0R7���X���u��ƈ���0bٯ�����߮��f{
êQ},0:�rf�D6)`�R�ua�ǃHbK�^J	+���lQ���e��/e�s��C�$�9�O�Z��,4Y�q/-.i���C�w�L@ p&f�X� ׫X�g4���d���o/���a��囶[βqR�&)?m��hyU~UL[e�?V=k�Zb�����&||cj��J�z'��B@��l�*���à{�Wi��z7��N0\t�MI=Mkm�M��=T�H6���S�^�Ҏ�]�	�΄~����+[�_M��)�-"!�6�#����=8X��6�a	�J߰��S2�i���Սe�䇊�_�(h����n�����u���]L�.Чl,�=F�U���N�D�F�R�XR����EPU�N���ِX�����q��g݄�RW��1�kA��x;w�a���g��jܹ�lGl��o��/,��b����ylE�̙f����JI��Y쇖P{ �ёYb;O�P�m��!L���Ө5��2O �ҡ
q����&1��b��*n��6�`��>B�s�I�a��C�`��:��CE7�[/m8����B����+�)]��ENu��(J�l2�và���X����X��Ҁ�,�}���Iȷ����V��WV/���34�,��s�j����E�Rj���;��e��SV�Z��Qwl�)����F<6.��h��N��i���{�s�ov�),Ο���k
�Gf!���R߫��`��X��G@�������se�t-���>��(��XǏ
�W���� |"]���?��Oy��9��uz��\�M��j��m�յ��z����/�B1ii��*�Bs�K1+��In��\1{��j��k�Ȟ�L9��|��N�-�<�v���֬�BY�r���Ex�'dLd�jH��Va0��bD$T�^]�6g���Z���w "x"VW�;���������;t�غȿ��)]� ��C�zii2D�29�V2������uۏ��.���W��J�17(*�!�v�&�m u�0�O�-a�?���, Jle`�1:wFХ#>�YKu�Qޜ�Xk32t��p�h<��K��h����y�B��s^� "���o�\lh+���ʵ�+c��Xu�W.��KK�/���ڵw��*!l�%#H��@��g��E�bB(,D���,��}�_*:�aB��[�k�Y�����U�쉤�R��H{�<d��?�-�->/2Kf��-@޲ϳ)�Or�+E]���<�=H�+�iRŎd�B�ٰ�|нi��c�g����o1p8D�t����x��P���"7�
�'T��L�͋W��`Cd��[�ް:X�����'V��~�sH$�|��A��d9�zP��z�� ��m�P�(Ac�D�M�;�!� ��!��[��=Ge���	q��V<>��G*<�J�\[�����rȞdg�"{��W��U$y��t�"�겐{�+k�X��+;���i���Su{�~
�$�i|l�" �i�j�=G�����{C3�9������p
.��	� �BpT��o?�i/i��'M3|��?��T��"�L�:%Ö�R�1s�\�����!�mxh.Wkw��aJD_���.i^jg�ۀmUS�$=��Y(�rE;�?c)�����OS$�cS���Mҟ;6v�U§���x�.��&�cx�ix����U��i�������;}q7��`}�J��u�>�[3;t?S1�gw�D�ж�a�#V��i�#�����KM!IY_�R4�K�r�U����hݞ�\孲�������p�5�И��*���q�e#���ĵ�vE=[stcA0�M�0��)��t[���*뇟�����)�������E�.+�L�_�W=��B{P�V\�v	B9��6�����I����
D���.�c �P%���N��ݲ6Kaj8P��=�S�1��49��e���R8�r:���.�qkpcuR�>��{���VJ*�Q=b1���Y��Z}��|afW�?sR�m���_t��Z��bT~�o�׎]Dj��b�J��#t�y:$���`B�����6*��S� B�HI�1�?�7���>��ECa`�4*\�\')Z���d ����Mh�c���!�����Y��W�7c[� ��Oi�,�)����
VĤM�dٵ�w���9m�1!��AF`�I����v�Y1w��g�i\�:�	����+M�)�B&�~�u�zK0-�^�tk.�~�g0��?᝟��i��
�vn�)�������՛ЂQb{��pI�	@�5V�&&r��?�#y
!@���f���L��!�qs�,]^f"�{\�J�f �`��ڢ�A%+0!���}��d�=�_���CkY��!B�p%�_�q��G~�~���l��px�%'A�t9Nѷۼ��IM��Fهp�',����p���	�Y������H�^����zٗ��q��D[=�¢G	j9ġiGw�OQ����D���e1�+��G��Ve����rr�D��N�("��A���������:rc�a���F,�g�r�Ϋ�I����7E���l)��KG@3�ܡ٢{�Q�k~{��d��]���Fh�<VY½��+b�;��
����/|D��v�6qU��NmA�w�����e��1|��~�߯&�g_
�fܡU�bGcq���(��hg�����������Ĭ�=�;��k�v��/�dT;���^��|��+�A7�	5�Y�xlm�u�:�B��R>�~e P@��>)��m�·�i
�|&/�O7�;(�D��To;_3V��`U;�I=r�T�/��ޮ
C�so�s��܉��!i�A������8����\�i�����@G��rǱ��3`JQ2"��oO����zAQE��nVQ|
�m?@$�Lpq��^���zA�ߛ��W��~p�O(�y�D�_�;��ٿ,�u��7#�;�$�Z߮�R������&ץKG��
���m�h���Hu_�	��W4�F	惝:hd;����7�d��pi�����;�#���i�2,][�>�\�i�B�#�_�~b���՚/4����h���!T���6O2Y&��T��>�I����ڶ[�qB]����&"����|�l���?�"��+�؂o����M�c(�ۮLu���'�M-�t��W՝'Y�lщ���)1�N~ B���;؛Z9��.��߻?K l��=/,���΍
C����H^�}�yX�v}�t&���Q�!��|�H���9db~#v�{K	H����x����q��*B	Ͼ-d�����2�W���	�rn�0�p���vm�|:�r\??��3�#8�dm��9C�8 ySds�5��}V��b$p�a��g����e-������=C�� Ϭ�7�v{�Rdͧ�Yu�z\��y�Q"�j�.L�<��:h#�>�u��u���߷���8�|j"�\�3��I
N���"렏�TPC"d9��+�Ak�M
�����Z����Q�f�c�Q6f;������.3T�cc��Y�sb�0�;�#�2$Ua���I���Q�
K_>\[H���K|��1� ��S�T��d&�ɫ����.�O�n4m�nB>��$�Bj�J�8���Z�ʣ4����K޸�����+,�.JYXnNp}P�+��`+��*x(i=:I�.)��&s1=�.���)�R�j ͥ��˵��YB�5��k�a1LX~�}GA�a�����W&PA����I��>*H���q(/���vnځ2�F_U��5������7�۝����m�v$j��(I�P'/f�r�&b[�*7��娯�R��动�BfE�K������L��4��lm?F�pg� ,�I5B�����b����0CL�v���a�D��pu����(��Wg,Y�
=��[����%�r�7��C�J��k琉�L��2uB��9<�Y����&�`�`�I�D7�G~�y������ǙK{��u����2q�S�Gϓ�j��6�Hg,��d�'Mn���ߍ�G�Y͆�Y9�Cܺ���y��A�'t�r�V��AT����E��q`V��V���*`e��x��
H�b{B��▅�u��r��8&���a<x���2����YF�S�׊
�)8�,'#ѭ�1ױ��=�JQ��[��Һ�#N���:�����+ڞ�Z�?���4��8��r��v���7��}q�o�s�R�J�0����,5CU�+�[�!��lT�6�-�bߥ��5��� ��q�)�_�z�=��݂ê���Ae�	�Ǘ���.�H�_�K�n]��<q�r΀P�i| e�Z� 
�Y�g��X����r�O�=�����R�b}���Lɪ�F���!1n�9�y�wi08��	{
Y5pw�c��h���A����@���ٮY�}�O�EG?����Ju%t�7~>��菓QԂ���{H+���g���}l1I�!auc���%Κ�>�7{HVȪ#5�ᡲ�s	�
h���˞
�/#M4�W4a9PZ�]�(Y9�Ш��Gp0 VJPWm�P�h����.#X�z��ԧ��ǣ�,]u�l��&����
�D����1���1�ŧ�<���w�gvo�sH3�45�j��Hځ�9X�1�j�'{�9�c��J�vQF8Y�-�D���ߣXo��"fk	��I���6-	�I[ ����.��]�*����%=7������ڂ/����������%2����I�U�8�e��m ��+��%�q�iU�X��%a��Fi S�Z�43I1o�%�D�$V��	��yr�K�Y�B�fǒF�egS�0�ai�����8�;��o"�Ҽ��B������N�@����j��a-�[��ޤ�6q����dJ�/��bE�'�68/���+���Bҍ���)X��^�u<R�d3���ϟ�B2���!�H`>`�*�P@� �j'���U�ͥ5#���`��=R"�\I������Є� O���ɘ�Z9fh�;���5�uףԿ�G�Q�:t�c���M)�>���Z����j���{̉��a�8���2����왵��*3���G3B�Z$p
;��G��Ϟ	<j>T���C��"���a`w��#m�{��k��3�^K�tب�=75�p��-H�e˙ڏ��?��g�{�@�Ǜ�E���@c���E��/:��E�� D��w�M&�D��'���.�=�����2�l��v��1���������J�ih����ɶW^�	��V���qi�7�跠��_�gcՉ�}]�Bl{��R|�5�G�Mow����~�Qs��2�J}��f
�B��?"я�-~��३��0�N��2��'��߮.m�>/e{��(��յ"(:P]��٣0�u������)�<\�Z�%2�b�{%�ew'8��>X6*��+��$j��PI��鷍!�Pxg�����rCy�*?yY���]�ʞ�|	�f���~�����; �Β���������RI��D���P8L��i�r<�]���觵�E䶫��Ei��mF�+H��n�b�X���:�7;�]�c��/��ٜ/A14:�o�$88P��2��y�"��w��&Y,2d�H��|/k�(�4���=۩/~t��>��F��wKRD|+���<�)��Εߤ��Y8Ζ���)��N�{�W:�Y����q�"U�V�e�����c}��"W��ܧe4х�1�r5r�63~�����`-C�c-͂��%��,t�PǏ�AR������gq�鷚q�)"@!E��Ab��7~X3�͟�^B p���.�����73����}�*��G� z\U$ٔ�w�X顭�^A��()�3�Fk�J-5�kY�������:Dh�_B3��d��?F�0ri�v������5=_苼�w>������J�G�JC��]�5�7��c�(���PF�Z]����T��h�J8�2�J��>�������-��wס[�{����Т��uc�|�|
�L[4[��\r��7Dfԝ�N��z���D=ony˴�4�V����*�v�Rc,~BI!I��9'�fs#f]��[rj���B=�'���ˉX�tx׻rt��U��^1����4�F�G�a�fHS`��׾�"@����3��&)�@����
Ϸ��x�������*C��z��d7P%�vei7+?���������h=��j�H�y+i?�^���^ɖ���E��_\vs/'B�_�aѯ���H63L��)��<�~���G��*d�_����T�˗������ϴ=��*s�Ag\f�j�����D�t��x��SU�G�^~���I1q��Љ� �-�%��k��.�ޱ�U�	�Zf]N��y�B�
Oe����V�ZPc'����T��N4�^w+���N
��U" �JF��u�&�]"�uwQb�He�q��|�.E��������e�����$ ��f�A�	�SS�=x�
U��g�eկ9����E�z�)��Y����L�6�������{+b�K@���N�;�@LN1���fKouј�/X���9�$oﶚ'QwEHH�<�L�����҉DEK6�1�i$�(%eKr@�!S��O��:�H� ��{\����3T�����	v
�ܺ�D\�u{���{q�^�Bm�#��U ]9��DM�/��������|�����U_�� {�ד��g���+�q_��U�<����!�cO�n���2�w��5�z�+3�C�$���K��
���7 !lW��^/SDuϢ�{Qˌ)~���.�ҭ��-R�^�B-{6�:���.�דl��08�Y��:��|F�[ŗ��ba�� F���.�֞pB�e~�C=�����c��c�1Ù$�ᰀ����B����������XJ7f�yoH�[X:���I��Z���n�����ţia`� ��T�r�a��4����RZ��\1�w��A�+R��ʄ�ȌA&�Ը�@�%-M�ͱ�2�)�|ǰH��*|S��~'\Oa�1�!�&Xͦ6J�r��;���Ƹ��_9��F�ˊU���>�=�h+WQ|�|E�0��8%��L��L�X^)��2��(sՃ�y·=,;."	��l��`0�ʆ"+ @ߨ��A$b>�γ�0iI��&�G�ݱ�J���q��(��q��шE=�;�;� ���7'�g[ޒӁ������޴0{r%fF3E�bBT���C�bq|��'4�l���K�_I�N�C��?�������+��e���	�`��)%���|��"z��"ET��#�<��/v��\F���mt�GpO�G��h���n��\�w�m�!�^�<ʺm�:�$���2�4��AygH�*�)��{�,�����Gѽ�8���4D�2�33�Ԓ�Oi�Me�h��I&ₜ��4��}$�ٌ��A(�T��^%!��D[���l��N�Q?��g��@��4�"�S)���o�d0{�UPsI�E!2:������kq8ꋜ��5_���4[z�0�s����}+�NAt41�:��RF�A(`}
��8���
иwͪ�`=����^��@V�u�����&!� e������(�&�f��N̓X��F��NڌN����Ҙ?�i��ܢ�?>�}�.�����U�����P/bn,�����u<�XB1�K��,:�б���������27#��pKDA.�]ާ��c�X�O���I�w�u[2V�T�S����z1�\�τ�=�#�}{2�[6w!)U;2Ƅfws>�����ǆi%#�,aJ芤�&�Z�T�h�[!�K�b�������O�2¿SR�nN�9������B�Pݾ.2�.�Z��'�Y��d������Ec��! �Gf�eN6f;�#������Pw��5�
�F�����7�t��IN�sT��s�wPCa�aT�h�E�<�s�� Q�dlZw���@�bN�i�ê��hֿ@<3��z;Ks�������4%�(/��ٔ7a��z��/8y|`ӹ"�f�k���C�q��j���A�G0�u �<�0xq�hmŪ���Xr�A���Όl�S]���)�����Ld[��.
P��&���*�#�Qf5��R�R�@9� �7 )W����ZG���=���	\�E���Ï�I�n���A}Ȏ8FHV���zg+|�i�佧i�@`mL@�Ȋ��J�K{� ��{/H�~dv����;j��C�ƎY����z�l�v0/ ������I�����zt�:I��1]�"�Z�L$}����7%iDCQIau�:���6@O="�b7v�jiGZ.i��sxe���E�� ��e2C��
�Y�i�+rt�ƝgOD�i� Q��hJ��:	����ڎݶ3d~p�7��1qjݾ�Gܢ�,��2���昅���@#��3%D���~��i�C{s7ERFt�$h�ݐ�����_��a�a�g���Ԓ"!�(��x�uTx���O��Fǆ&�)�w�.Rx��z
�IH���lp~~t�@�,���Y�(�0��^���<�	�� ������rxp[����Cρu� [�,l�:���G��C�ƯL����
f�TTME-zjN|:3�
�hF	�Hu�����TX�k~�pᐜ�kE<F��I��/B���d5᧰�sh��'Dc�ZkW�X���� ��D���SÌ>�x�� //B]�O�;׻���e��*ֈ!�v�"����ej��D�؁q]q�/G�,ʓwk]]����M-}y�V0�_����g���^(vP%"�t��4`��
�qu�Ô{�h*U�/��Ƒ�/[���Kr�%Cz��l
c�:�`3<�o=��"�ַ65�F ��:4S�o#&����y� �w�7��G�k8���w��S�3Ȓ���}"���6B�����`΢�px�d��,���_�L�8(��*�c+�����]4}��6�4�h�Z�g����0�8W�E��8�ԗ��{�aW1F�0�H|��1O� 9�e�xG���Q謫��FM�YDdY��ٌ;��^�$�agi偢F��+�>���7\�4�!��6���SZK)bo�ܾo��~	�։�J���$E�7)��ը�5 ݓ����5�?G�����>�&N�Qi�pQ�/cܹ(���(����9?�������+���R� ��D�� R 	,���9�(�w���{v�.�x�q���M^��b)[D�5 "Q�=�.�5;�+&�߸��c���Ǚ�R���|����3�5�,6hk�� �9
m�K���㝲q��ɂN.��
V��eҋ�b��ѧ�)V`�G�{���V�$���8N�;W���Ć�m��\�3s�8��p<.��nn���D�n�z|�*VqY`�Tfy�7S�&W�+{Yn(����w��G���H�A&����i��-:��N��d�^��"�ƛ�}A�o�XY���l���n�}�G7�p�H�hK�Oì�RoL�%p�+��iÑJk[� ���]��j�8�_H�?���%I��|W���r䥟�xIҰ�ϥ<$��?��� �H��0�H$a��ؿM	��s�>ݶ* �����WA�+�jI���\v*w�xN�?.}מm1�����!���8�g�Pe���5�_�_*w�B�������{�9�E ����m#�gnn([�z��l��1R=Z��������X��3�p��`�������`c]S��%�v-z���s��c
��dl�o�'q]ǹڊp�MW%Ӟ�Rڗ��U%:	�ל���(��%�Ya���s�2�L��U���Z(mE40��C�{9tOk��2�Hb8��KO4�Q�.o��w��@�{�_ĩ�3���l�ՓV'vzi�yq�0�H�qa
Ͳ��6g9�R[dQ�yNZb�հo�ޓB7ˆ��C������L��Z<\	�v��i5��&�6쾧u���i~�1��>�B�Ghr��G�.N��ΡZ�yV^"ɛ����p �Sg�2�P���*G0'�4��'��P�U?ϛ��9�פ�z������n�P�fRs9":Y'�qPQp
���lڀY�P������ƭ� �U����s�wP11n#5JT Mm�1_6G��L-HQ�~=��H�������6���,'ϰdm	0Lލ���}���t�X4������� �b@�aa��AX0��ߛ���&���~� ���|��*G��ձF�Lԏ� Nx`-T�J��ߡ��_�VGd�/��]"�3�#`�y�`�ߎ���N!Adf��dB-�	X.!PMYs�"��j�
�jѣ�򓠇cj���y��JR#>��8u?I���\��-QB%�@�&��m8��#��o|	L#���W�o��b���?D�l�j��/�^����M~X]�o$����(�[c�|���鵆 �:��#� sEWWb�s��%� ��j_<�_���I�B�!��P���>?�.��{I+e�Lvwt�燆����5�T�	Bt�2Y��*�|b�^=���y{X'V��߈�]To��[�A�߃!J�˛�}���]��3��{;G�u�_�������p��*��ia��s���e��N?0i��1[�0|��8�/t�K�ݵ��/�-<:�ġӼ�Bku�?���;�u���I�c�qC��<Ԑ�JQ�y�P^��D���������}��LNV�ל����WJq&�oBXT5B�f-��Y����>&-;���Qq��7ʭE�*�i�h���5g..����a��n9%�[��)�?*�Y�3�<�]����0/�]΋71��j$��ļ���'�}�ȷ\1k�.��3. E;Q��<�?2a��j��a�#��+Z�� -��uT���kEGj���Z�\ˠ�U �� ���pI��N�b5�6+�(�\��61#>#.��H����u��*�|O����Z�3�� ����o�j��e�d��
����W�����v�!{Vs&h�4���W�2�/���BgɮNʮ�|뺘T���@�Qg��Y�T�	�/���}h�g�$�CX��{ȷl��_?y�"N�qpkQ�Ey�c<17�a^3o�O�m�ߖ"֣Ϳ'�o&ճ\�-F���p,ơ ��_ ?`�������Q��ʻec�5'SW�v���(7�jQ
^/����15#:kV;g��Y��\�6����賕Y>(�eDHiS��V�}�������wk"��&h�aH9V�����K�^�����;k+S�K�vߨ�		"F6�x�����k��q�:,����H1{y��$iN6įPm��L ?	��|d��m)_:��(M-���KY~���C:,�/G��?p��Aj��J���r=����w��Uo�a �>Y�f)�K7"��O��3�+"�>c��g#ʁl{鐡���nKa��R2o�P�Ø�y��yo�Z9bE�;�\_���7��u��cY����/CE*�B&�,D��g��ʘ&;��#����D�y,T�"��_���J?>۷��j��#[/.�K[/8k�3&��1�X�y�J�mۯ3QG꺼��������Q&)�� F��ׄ`p��Cw4�s�u;�l�{�+6�sr��n?����Ɍ������ސ�ւ�`c)a��^�_��&�'�?ҽ���@^���=�Ŏ�q#��b����,��;�~��-=��c��V��g2y����Y�i>�oj[@�䱈J��[��x����bDf&�(\p9�s�z\n���{��W�����r�B��׈��`�#�<b�5_,4���~�7�
�Suh(s_����Sq��ғe^n����k�bK[�5o}�w9化��g������;?�	�J7w��h���5��k�U���e�����D�ZvF�$ҡ�9���:=6!�c��U3���b�:�[��c+j�,(�׸I���\�W��|ǉ;}՛޴�3m��Tb��x�w�"VWv>J��u0U�X�?�� �&tU
7���Y=Hq��U�?`aWv��.��"9�=�e5r-��	�f?�wʿ^�#����
�j���������0��� �n�E7�?�.�Rt�"�F��U�Y	�X��}�Q��jB�҂�DA�{��/z2�./軖yCE80������?Z��
�[ޏ�C�4�+Q`��+{���s%j<�^t E�Tݦ�����ŝ_
����{Ѹ�F@;��.�zom�� /N�eW�Y�%	A�RcB�C����)�����\~�����V`��rx�x���j�����}�%�e�8��y���r>�g�,e2���N��)�;Sxf[}!��<8��tw��cy�=�*�(:��܋9Q���I����bf?>1VW\h�k�Bߢt�M [	�̉�"7N��N�l0�w��e��&���[���2�ߝ�r����9�*���W'���|�5��vy�Z4眩�?֑ס��Ҵ����L}R�e��,��i�:>��oʓ�p���bwJ�"�|�ۦi��_�i*�@����x{s)[��T.���暎���+��+�ñ�c*��mE-�䷣�L~Z0���K�U�'���6��<L����?���f$'��������]���}�Ƒp���3���;� �M���*OhtK�ϡ��@@�ӹ�p��&����$=��ύ@�#�ߌ���w�18Pc�_�8�'��%��\ᎂÙE���cq�x�l[8���VB�h@��m�3bޅ�by��4�R�Ba�@���27}v.��^�;������������M|Q��e£&���)fIɡ_3��/��d/~��{����%D���d�N�;�Ve�o
,ZS��(��?󖕉�a?+��5@i_�R��
�P&Dw���y)�ջr�	6��y��8��Q���7l��3M�,�Ыj?���&���'n�=�5����l�T���~Q�UNo�"Ҙl��k���W�uЁ�So# E�g!\�Y������6p������7�6�虂n4�����[�W�'U�x�����N��'�s3Ԁ4�9�yK�|e�o�Q������~�H�,�?YO�H��p:�������h=��N@p�R��މ
n8��G@�gL3O�_������-2a����r��0�������T�1�����aõ��f������M��J:�=�@�x�&���B�?%��ż��/#��2Tʅ똒+В� +m�i����v��З�,���	..x��R�l�:����C'�H�I�%��(,��hx<y��O��X��qx3��UȬ�@p��M2h� �n}n�pO�@R�eZ�~=�O��#�?���+��"��^\�S�|
��c������!�K$I��>�"�p�1�������?Z�u0OM�1�M�C ���k�A��?0����1p�3�{#tz�Ǌ��%��NW��׼E�}
T��m>X8� u3�i���e�>}"��r�s�g��h,|�/�����Xj	ڏ�?!e��: �]C�B�K�.�s`�C�b��j12c�d	�n j��U�럵��<wNxX��,�/�Cd.H
O������{8�HO*/��7f6'^W@T��A[ �XW^R��.���u;����ʽ���9B>if�����|�V(��k�h}S�H6��q�_�8
����g��ǥ�)4�-ḽ�KO�v���~�4�4��ދ;oj����6�rHIP���װuhNqr{Tp�ks�����JXJ�/�L?Zo%b���@_�Gy�4�NU��JAD���e�Iy��ŀa��b�|��=��/~΁q�1KH"m�$m����ՌY���wut)�����%q����C	Ҏ�q�3-eqH� )D�ˠ	�m���iӕ���j�r0�˽�&؃�]Ԥ�%ZǇ���4b��X}ra��r0Qbn1�5IGV��{V�Ӛ���c��j�=1W2{�&:���=[��M���4h.*KE���y(�9�tB�>Zru�27y'꾟��V���"�x�QР�+)������[�Vm���ݗ%�--�#��������+���G�ei3�&���Ty�x?�'��$�ef���x�Eř�1G�;�jq�1��]����"�[.9��8��xC���)˭�ö��7��_����Q���c6�y���Qν�蕓�ڳT']R �/��v�b��xN��觸iC��N2��[?�_��(JӉ+~宰c3ϫ�r�;��nsc71Ó��r��%}��~���у��9�e;9��H�k�)#��%�sq���__ũȬ'0޽�Q�*�>��w?*���+��kD�����f~鴄p���sX��?%b,b������0����)��@ݳ�����
�h�7�z�R:�T��c=�t�N�W�mCh"�l�n�j���8f%��7$Y�(�of�Sa����!�`5�-��LՏ�O��+㇍:��K�s�8����'#1n�m;�بR�F��9[��K"*��w�Z�e�b*�6��A�u�mg.J���W�i�+h���6㦂uZ�S��¾w�,θq��ܷ�V�i�,��k��`��ˊ�G��L\^�a��ѩq'�QK��0�Ȋw 1k��o�FP}Q�'ּ��a�ƌ��+wcZ�� ��t_)��X<�@�̰(�����������1�Ci�{�� �PV�qn�6{8&EeKt���0� #��Ĺ4 ve^ӌ��p?�=C73���&������i8����[R��L�פ��]{_I�s`��&� OY)� [�����TR�{�+yS%�!��O������ƅ �w�1eX�;c�$@�F���Ͼ@��])�鎯��I������Mі�����m#͈7 (0zS�jͯLik0��D��V��A+VB�T�0�a�)Șf��fZ����*�;���C�$�L���X��O�e	�*�?�ҝ�+U%�8E�RU�~Nh�E/[?�ٵn��q8��4_%Muӷ��s����<g��Yt��8?aXƦB \g5����ĸ]�Y����M7��}�	L�_��B��c�Y"+��F�z�Z�f�`J~��d�I��e2�)����gX�������#��\?��ơ���mK��O��� ��x�o�-	r���sA��^�]'����E�dV�
"k߫9��b����Uh��K�~$/ݧ3�C�*�O�	\�[/�θ�a:n�N�im-h��C�+:�H1�n�r�è�<��%�ks #��w5Y����5���jD����&?U�ӆ��ܫw~��:0v�c�Xs���XzU ��,6E��������@�|'�c����rђ�K~�����}x����Ɉ�%Q��1{��{�cՖ-�A�����R�g�^~�&dg����g��7ny�_9s����R9��o�&E�=7qag$��l2Rܣ�Q�uFD�p�){
�0����}9��[۠O�p'�~i#��+�ԖA_�O��-��#��Y��nh����ؤM��M�
��3��q 6�կ����'�6<0�9�����Q<h�w�� ��x���'����D�2�LiQH�i�,�2�7�\WuDﭻ��}����LE����M�K�/���צ,��I,U�*i�ԯ�+(	�X�p�i�����K���	}Ctr3$[wW|��_�������{�+ְ���d�i#)�,��� ��|���=����∿#�{�Vz{�8��x�~d��L?xl��f�к�B-ZPg�i�m����s��t�����������_i��ur%�X�V��	��H�UhK�)�����z*j��<�&�t`%;F��JD�x�H�Џs�|��=a��0�N���³i�MR�q[�je�4XX��Q�v�2��"9v5`�\D�ssz�!�4��	��oeU'IG��K~�Gv�Y[8X���?��]�7�e�PdP{Hр�ǟ�l�����y�C_=1V1{M���UGڂ[,fɓh۞��CN^8zIy��>����;fAE�l ���ዱ~���Â��4ݜ7=�� �.�JNbϼ�������Ҝ����,�7�es��/�l(����p�T���AӨ"T�'�N�"�5���v
l���pv���0���8�Ab���W� k����a�<���C,%��W#���֘����w���3�`��Y@D�{����y��-���gH+ppΫ�v�65"��Am�Ǽ��	*e}���a��/��/Q�oS��LΜ2��]�[����?tHl_�LĨuT1���_{�z��K����L\�G݀x��/���做�"�$�dcڲ�O�K�xe��������S�E[t�Ƭ��_���b���R��ZX�Y��L_�?��V��x&E}*������!���#[;�F��Q��^�Mcv�Z�U�FA�vK\�V�6z�!��7�h��1�Q;���Cka� 7Ge��d�4�jGP��+2�K~��Eu*��� Hҁ�O�e����(�����x�8V]�|'����?��$u@���q`���F���]�,G?sMv~q̎�������K����[��S(衾�㵟II�&��+�|,<�0ʪ<�_֣^y (4C}O ϖ��C�8�C���gt^���h`��f���ۆx��pu1,��ih�jZ�Țn��B@��G�<�(���m�e�D����@�Y$w��yZ ��7�)�N�6SE���E}�����g������f�O�o�+T��0B�,3v؟��3O���ހ��o�RJN��)�@��F�H�%<^M�!�asW��Z���C̋cP�]7!\}'/����~$	^f:�Y�f�ݻFqe ��n�F	p}.�ᴈh3����	M��aE��!
��E�S�O-�DQ�&H�U�S�}|�s�^	��g�����'3�ʄ�D�:Rj�1�iܴ��.��%b%1��p)B*�� 2��j��.L�Œ����V�,��,Д��|�V<}8ۭ���أ�Ţ��D����♪ZD4̅h�	�k��μ�����|^IF홓�S��t�	Qd�p�k+��S3UR���n��mr�n �q�a�t�0�����U:y�~�JB׵�5����v�J%��a�q�0��-�.u� j�s;�~�T��S�O��b*��]?���.��]���	���s���u9�p�ĥ}�tl396�I�$��A_�-���-���yYڳ�]��3�o��@���a�y:ʻP[���g$&	/�k��gl.��F&�����z�ڼ��	;�^���[~���O�Q��h�
�w��w8�ps��� /_����b[_8���k��++8��,��~�[���&���c�1J����)h���f�p.p���#�3����0hQ��\$Hr��`�`"	�\	ę�T��̧�~�����F���!�^jя\�<ˠ�	/�L�գjl>Ъ�="��D��J�5��*يo �˔�3HsN�`��"+�!^H�N��Ԅ�(�hSXǾ�sV9�tT#�d�%{�=�\�:��L�ѶJ�y0iv�����M�?���-N����ԄZ�g�y�e*�M�R��R(�a}g�4-h�A���,��iG����:N�p�2 3��<�\E���I��<+� �C/��h�퀣�a��>e���ӣU��P�'�4�t�������mP��Dݨx�1SS��8#��q��(��W�S�3��П����eD�W�Ԓ��^��e��N�@�"f|���k���.�0��tm�;P�]�Ϳ�Ԝr�6�[5�����a�_g�֜&jSt�;PŨN�wN׆���I��ȃ=r�!{��E)*Co�,M��?,�I�q�⋾�	�e�k^��Ds�fk|QZ+���7,��3�%t���Zď��ϯ5��B˃	�e�߃*���&�����e���I2���J?�r</o&'�.��V^;����0�8m��64�=_��U�"�Z3�Ξ�`��l���+x|���-���xOuH�z�W����/(��.7���l-�e��*
T����Ơ������~��JT
#�>~��~F
���T�d@/(��W8�6�0�5[�� ��I!�g��(H��d�zb��k~���_���N
�z�yy�oQ2�mǓ����7`�r��<�Bw=?RC�"$�rv_c���shQ�NI�U#��^O����I�֬V��x�ey�B�_�$i�*�A|3ol���\/0%S3�z��"Tzd���Sr[KX���@�s?12>]�0�#GGR����Ls��GxuV�<�*ϼ�}�I�w ���TObd�hPoh�]RQcJ��]�����;��n�Y9�j�~���@�/���+P������1]����8� ����2㍴�86F�r��"'`�BŹ`,^)<�p�*�A$�gX6l��U�u~92���<[	i�XUV���{��|��	"�m��aD6��t$n�פ����{y��v�y�,��ߵ����ҝ��$ň�*�}��Gk��+����q
�--˛����P�+�MF�(s멬DL�/D�Փ��ٳD�|��x�bp��n%O&����qBD���ք4bl����Yšx���)�w���&;z�NψaP�GW�� ���d%g�R:ǈF&��I��"�4#1�tU��-�9ynI�X|��v�A��t�Ʊ���Q��K������Z>��|�$�\ja�7��wH�s� �/J<�܇���ǎ@,�ƟݺT��\|�P�%���У�~F[U��@_��钑� �5C~�Ã�R
r�1��Ҝw��H�$4�J�	�tm���5M��]c'�no%��/����C�VC�/�V{d1xAg�$ы?�r/�n���h�QȊ���B��ٳT���TP��N!��{^��w�R&A~��ٗ(I��x���"���&�-v�
�ŗy��<�؟�QD��{�i���a���7�N�|n��|���C3H�ْ|������
��o��u�
k��п�����t�+���`u:m�랗fb��.�1��:��L� �6C��S��[�[�h_]ClG��S�Ѝ2@Io���2�*6�W���pBͩp�䕲0km�űx����ֹ�9�N�ݍAxm���� ����#�3_���d L����+�!m��&t8�jw�q��7�T�X�$'O�h�ɚ�ץ,�ݡ�z�4.��sD�Ĉx f��]7&`lY�~r�+ס$�1��ėOX�7�	զ���X�j
��s�^�ŀ���d����~$Gx!`���Q������Ay��Rz퐫]G���捁�k�z�d7��b�	�Y�go�"��ˢ7���ޕ�y�,wc��J��?@�V�O���~�t�a񖁛X.���ʇ�V$�
��i"�3�������7�>��م�3�0g�YG7+ש��<����j��mCB���$�~�Ծ�"s79������7��ۚ�V���};S�S���.2��lQ���`_�s��n���)����*M�}�8-{���[*L9�
��5ϻ>�z�w���Ӑ�x�4�,7w���T���dV� 8@�Y���3�?Y���a�g�~�9���j#,�n����[[����1��\�s�ڌ�q�c�8o���͗�����Y����L��x��3I�!׏)�LSv)E�E��Ԗi@��H�*8���VT�B��\�!�j}�=|�����]�!��M�4�t�P�K}�j�'�R�c i�ޡp�5��)=��vo:��s��b"�o�6��rJi(C�;�Ї��W��B����Ǔ^��������CH+�'Ky�����N�Fم��i!kf�kݎ��îKc�WR�N��W��5j�{c@s��r�V%��Az�ܾk�4A?�m,k�	D�������\�E��GJ�L�䄷�#�"�L���`f����l^��[?��ݚ�nH饠�Km�+Q�*�,"c���I�O7�&�!ڡ�̦��ا�he}�c���O~����(�D�Qֻ�����]�w�
�U`�Nq>�ԱѶ�<�֍m�`��h6�e�]d�hIX�Q����{Vt�}�Ly��r�Mh�6s�H{����id�a9�kB	�-DU���K��8�����;ٿ��AL�5�br�Q�Ds	~<�����Q��`���K*��j˔ꛪ:�ΑR�?�2`n\��i�ԁ �:z����4��������_;����cq�5��G���6��~O�Yoe�㩨�Yv,^es�7c7�%��xvz)�@t�/�VzD]�5=xA��W{]�m��JW"�W��p�x���6��~r+<��^c4e��#��v��1$jQa�03��B߃�d���ţ�9���3 �O���>Øz�H�]��hK�����g��S��Tr���HE�q�
y�+�ʂF���ϤI�OT
�����#���7F�l!�k�XS���|1�7Bw4@bq�	���y��C���� Jf��M��0�UH iy���U6�k�t�>5��m~�����P�������F�I�8b�C�CN�KI��n~7�I�9�7�E���k!'�i
���������<�+�N��	�CL���5��h#&�����=�.[U~��� �]#����ٲ�@�OR5��ŸJ.J,�j�J#����ʐ�K�c�T��CW��������r(��Z����բ`�E��)���1�]�wrJ�t�UO�V��̶	MzB.�Rz	�lB~�\�j� ��S�羄�:�q=������^vX��z����V��D���&������U�������w�rt{�m��i����^��vCv�=��MX��M�z�Ҳ�q�ўS�N��@�mM@�B�I���;,�vHJ��{�I���fC;>S�u��Qu��Q����5~�D����Fr����_g2Nl�!N�
C��}�sI z,�k����yi�(���~�?���qVf�
���3��g��Tc�aU#�7b������b�K��)�_ԏ�%&٭H�D��F��?�F���*r.�w�`����ˑ�-#�
�SɌ�m��ڮ�T�1�%�7\��f�\�l<��~����}�c�Y8�Ҁ&�����3?�Z�	a�3��rC�;���U���n8�4��lA����4t'i5���!�U�3c=��š8iY\��t��;q*%�U��MY9PW|�+��ۯS�	��يp�q����=�L�́ﱣ�H�uT���>D���^e�J��i��p���7���;���u��]�豗�J����ϩ�f�Y|��z�O���og�1���r���Q�q��0���Q��9����r窛�+�`�Y�fM����n�����:_Ƃ��_T�xc�q��3��&�#��i�/��B�\֏���[�]�T��m�#�h�MWn|kui�	�O���fI͚�1'	l����c��B�9�z��x�Ln��U��@�|�[4_�/q�!�P%��K�Drj�&�+�oj��؎V�)@�D)�u������͖���#L����m���̧�I�Ӗ���P�������]mF��!H6xW���0м,y�[��Q�o����@b���ˢa�Ŗ��t{�^��^�gB�r��ZLNZ�-��X�ω��2(�;��1��I�X�`�W��V����
�8�8���n=G����<l}��H���˩h�7�G��_u���ʲ�2#i=�^�X]�6x�
T�Kj�(�6���$}ډ-@�gk�z�Z�7 �fbޓ�5<���PC�����T�6qݟޝ���;[�Q�����h�W[��a(� �H�.&1��1>�-��</�3|�
�fy���g�f��ᵞ�G��k�9��
�3y��	�XP1�$�7��&�H!�:���~!�g^�SU���5��n��)v��@�k�U����M^����9AaJD;b�*�Ur��ߦ�c��?�U]��&y�S�P
��ntZ��]�3L����/ld@t�/��d(Sj>R�W-�qٚ����)8��僡-x7 F
�����fyI���1���B^�\�t!�?.��5y��$���
<,E�����6k^N�1�6���'��!	�٢��ǙT�d����;NU���ȇ�`�9aq�2%�e땪�.��:���Z��Wۤ%���ɗ��:t5L�KGydȞ���}NU21�:B|c���0\6s�%�����c8�M�~�n�}[Y�}w)f�jG@M������������I�v��Հ4d�H׊,u�)&��1�����r� ����k�]�0[g��~�K5�E> Ys�[�	�����z�| W�^1\{%5~su�3a�E��LK�:�J��Y��Z��e��l0G8F�d�#nR���� }���L��`;%ڬz|�T��K2���	��-Y�e8c�V�S 8���qr���1z��9��eD�x�x���j`;���!P��0��P�<)��n�q0ܽ�"{��'��CF�$�m(��	�%j?��ř��w����P�u�C\����&�%��Y��cm ;���2��w�)��]����r�CI\\��L@�vo�s�bג� ���([v�>��K(Y������4`t�M����0�鵳����K���%b����֘�����(!g�s^|%��������?ʇ��*-������TzT������qw��*\���G┓RM���$�%�>W`E�T��N�E=��Bc@��|��~[�B��*���4Ƣ�3H@!8	{�9���E&aZ�3�C�aUfb��P��Q�ߩ��j4QK��Q��zЄ��8���@h;F�)�Vs��7�'H�BXV����mS!5�=��)����29Xb=	K~A*��6k���BX<�`b�^��E��8��i���������e�d��-SU#Ԅ�ZJ����D�L�t�ǋ�_o�?�]
����߸�9.Q�aM�q�����Eތ��CQ��"3>"i�9Q��Ǳ�%���$RS��g]i�]�݈[p�e2Ow밥���>��D��cոL7��c�Q����,����D���_rf��wAC�8=Ӌ�����^�r1��s@���o����|*��q���T�܎��(lH�LCz��+�A��L3����+D��/���C�R}�[֊T��C]%�Q�&�w��Km�Z�t/����A",r����%�g��GY��jJ]�s�m������$s�	Z$ܱED�H�M�W=������zK��mmZ4Y����pւG n�$���hd�Lik��5�C����w���Ր��D�=q�N�X�Y\�+-�&�?��K:�\�1�tM�z����0t�� zʚ�E��0ӛQ��-�����/bB���3�/Uus���RWg�v��v����e�p�^��Pp�����~���<�ah��2�)��G�7�����g�T$���s�~M�$�С�������B��QtԜ�c2�u�٦e�xl�`w�a_��c'ƟƟxD����h#jڙbG�MP;��*?�9�'�O���
ڌ�b�N
�� ��0`���L����|���1(P�;��H"�q���3���:n�h�7��w��^��t�Hjf�$�a@0�u�T�2x�H������#e	��c�↡�����P*���?[�Iܿ�<O-c�`�);v�s�*2(�'�4�c@�v�q�[�S�� PR�5o=��1�zgt���K����E��4{׏�1���Q12F����k������z�pRGܑb�l���i�+> &�A}�h�?��ǡ@"u���l裊=�s�I��Bԫ��ЖE�8���73����� �>�8��<�u�d~�M��1�K��%Ȼr)�ܽA�2�b�����ǿƒ�I�s^)�P|7���m�5ǭ<(�^�,���Ez��YNSt�}���J��|�2e�W��np[�W
��3"D��-F����놆���Ć���nN���-߱t\�O�'_4��kuW��:�L��ӆ�f/u\��,�w�,�Ek�R5��{���	gb���9h�>��a��8���h����Z��RĝrO�Z�Л�`Nmm��3�al��.4!�$�B�e�#4f刘0g�i�Or�#w�*���#������Wڱ��4¥�8"�d��z��lv|�ʃB��CE�Ѐ6�.��'9�w\w����Ȉl������t�ѵ�jLѺ����a<�q�0�*i��|�1���InIw�^�?ﾚ��P�s>�ř%~a�zIk�H'�#>�-���{Z!t͡���R�U
䈫D������nԸ�%6:p�|D����M���Z��[np��]!Z>+���K,��ss�fe�{�0T�ւQR\��2�V]ZNF_����Ci�ڐ�h�{�#RWs��"�yO4Dv?+U#m�Ռ����@�Lh.�ˠ�f�$A{G:�R��,Pmf6��qd��$�R�V�ڣwh�'d�	�v���C_�ݓ�����޳a�qa�{�3��C*M=A�T��X.N��uk�m��8X?J�k-��u��5��9��S���$�^V���#Q
�\�ǌ�I�_
��!
����@�W�pU�"(�&����˙Ȋ�h ���g��g9{a�P#�	�>���{�������q�U����������UL5B&ƀ_�G5��m7B��l3u2~���p6C_���`>�|6���7C�8O�9E�i"^!�5i��μy[2"	��&O����h�w��?a�74=I3�`yd�[;�G���,�n���΋��-'A�U�|�D�n�$��_,�ĨŒM�����8@�3|"�_�yC�s���[�?�����g�H�zd%��x�Mu�D���(��t��6W�j�Z�o�<a!�	��+�Ԛ@]1�1X�!�s}-!B��ԃ��2꛷̕�I��;�ŝ���i*{��9�mG=��'�>?����*ޠ������]�+�U@����n~P�1�' �0^��_�W���Q����_��˭�6,�ƿ�� 6T9��b���p(H�G}f<Z!-�����&S������ζ�����Z��e-��1l�Ҿ�8�|�*�V�$�J�^�H  �,yL���ІYX�p�aAeM�"ᯧף�"��Ë��.ն<Җ������+���ha�����/�{t������iT3�ʊk�Ȱ�מ���"1�C9!����ό����c�J��c֌b��4�ZUӊ��3壛T��D�gP��D��h�/��s��#rE��F�35C%���H&ߡ�	D��3Oh���;�V�~L���^f{UhZ�5�6�6KP���,|f=��Ge��B�%�&�'�Д{��#�k8I�hr9A�G3�=f���	�M�EWH~��8�~M"��'��nRз2H� N��*��w�L�w���-���=k��>�؊֘\��T,7 ���
n[��Yz滩'J!=iB�L��H9�N5��vȪ�4�ً���sIz�+2N�I<�^���;���GG��t�+]�"\�f�o���;�p�����/26Z� �Vgܿ,��n�4�mPHïpA�tRk��4~#�PK4�:�R�����U����L��v=�tɶ-�F[��)�N��H\ЈXڀx��\f����n��X[��^<��R�R�'͊�!&xq*-�Ў�-�l ��6B{M�}N�*q0�7��t|�DzC��P��9����|����	�u���,�m$��ӣ4�m�8cTe�?G�경#���捯4�ւ��m�h<�ȼ���-A��3g�mr7�}� �S�)~��$ӑ�@�g�ƪՒ��>z���u,�P�@�|��8`���U�׶��tmߘ�o�KЛ�6��%נ/�x��#�(�*�ԥ��G:��*��sP�V'��D���	��B��������b �@��z'�0�!D�XY�'e�}Gj�X�.�-����|��A���# 0Ƚ�����\���i2?g(�%6*�D^�����H�ʹ�8k2�f��1��e5!�0o�=t @�ɫ�"<RjE:f�&..k}��� ��T鿖=
��\EB�d(-��tHW�@�����]b�K�����>��DU���!YB�F�O%O�b9|�*�1uf�/ݖ�s:J�r�[|��S��}e�2�Y>ڃq4�l�����Iȝ�~/�T�5��a��s,��=�+��M��ךʃ��9�fl�ߘ&�@�1:-�2����3pt�#�����U�}���t��T=�ia�����Q��'�� ܪ���� PF�W����d&j��S�Uhݎ����ϼ���ށ32�Fy��d���$������N>$���Y���<^k��E�>O&�7�-��cp1{����SyX�mq��P*��-u��:�DP�U:�:}��H:�S�zK�+�i�I2��z�<7G���"�����& ��
rH��	8�,ѥ9I*�=�v����W-;��qj�' G��τC����X/�| Gx ݴ��n�$�%�����ya�ꂹ<�
���/�\n��M��s�G9���柶�wک��D$������Lc��;<�1� �w#���i'��ӣɾ�p70w�Vb�D�ԃ�_�S���u��KK�\WA����JUhtOd	29���!����1��� <�CNz�.��6�S�
0	��w@�epQm��I��v�3=�X(�@�'���%���k�.�rH��wK$�E���;��A���L��;m�/2��;��
��Z--�:�����o�vS�tDl�E.J�`��*��;o�w&�'�/A؟�7M��j�*��ij�G������ d/J�p�E�y���c��b��t�RWQ6�a�or@�V����F���z��>�x�6��>�D�,8�?��נ�i��A���^��F�JJ�:J�0��|t�J��R,��3�E8�ҷԵ�?��on���nZ�nڒv� V �,px)����G�5�������Րh�	(g��C5iu3.�[����*�ŕ�Ѥ^��O^��tm9���䡾�3�b��Bd'>�N�W�����>zJ��%��%��7$b���ŋ(��7��X�H��/��V*����	NE�긧�V����m��C���$>�O����^6a#3^}0ͩ7���Ȩ��w~��r}�AtM	-X��Th�*r��2�~�q�y��(��mp��f��\�b�E9�|��$�g��j�ĺu�<@JM����f��:Jϥ��E��2�凛P9�6�#�[Kk�M�d'�
$�@LG���Oq�)C"�o����\�Gk{1k����vv�N�.�����!s:H��B&�wR2�'��F�S/�8�hA�o7�����j����nym�����VdTڎ�*7u���B��I�̺R]ް��!���D?���*���̡��zl��߬0����ڦ�A�_��I5ю�՚���(6�cR�m��]�̆�#����]��`�I��>A��(D7U��:BJqS��#�4��M���|�J�<mvW��p��D'�w�[٬4��L�;�.AkXUy�Y�����okA��X:�׀1���k�j�̐��i���u��&>|�#���6���":^���hW �b�Ƒݭ�A7��`�:�_&7��M��m;7E����^m{x=���/���	�(�C.�6/L�~8�߅'b� {R��_z��6�R��kJ�s����ŀoY;��z���U�!d0sڍ��W`�g�'s����9����D��+�G���Ǌnֵ��{�%��!2y�8��\��hG���T���Lf�xO�Z�yJ�믍���f�+��Di�T�a�]k׼�w��Ƙ��p�!� "�$D91�)���c&�eMY������ѥ�^��*���9b�]���z�f$��_�q.헜��w�*l�
䪨�T�j�?��