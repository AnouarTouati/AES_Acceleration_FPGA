��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P3K��$�?~������\͡��dk�⍥xm3T��8�׬����:@Ӻ�n~��6�*ݚ������a4�**�1'wO���?�N38W�'�T�u\�V$_c�2@T�'X��Њ��7x��\W���r��A��~�wz+?�a�,���VSq��vO����C��\�����'o��&�m�đ�3~f���P�?��p����G�~?&���W�cwK�\k`�.�M�w��:0��|��p:ϓH�m8�Z��^�Mr��6w��0�&D��S{fb�|(������y��fܯ�Gr�)�9�2_a�V���i�6艆in�}��샒P$��eh9?�wg$���9��c��'��Ce*/��@���(\����Q��4��ܮ�G�J�׷?��}�5Y"�nC�C��
��D�����,�0��+@$թ��y����� ���)h�
.�C0�22�U�C+��es�X�N]���h��waf�w� �����`���È�d�L��u�
�L��(�K!6�j͂������r��7�B%�="�I�Z�r]Rq(N����	�L.L�Md�;��Ve�4��98�~�ӉL��_�+�Y�<2Ve�^b���vv]Y
k�&�P�;G�+�(YÐ!	��� J�C;.Mg^-�5§bݾ��K/5�� ���cʑ�8	�i���V�m(�����<�H"W�{�/
܃���\D:��Pl�����N�zIA0�!s��/� ��3h��A~\v�1Lʢ�#�qvp�Dp� lѷ3�N� R�c��L�v��O�����n&,��p�'~L')ߠr1��!��M�ك�ϐ��s�@"TZ�
��� �`XS�8 �l����ox�ȹ�`�rb7�M�����Au*�>��d�7�_��Oх�>4�>��V O�B��1⫍`D�=�1׊�rE�h܊�;���,	����B�Ui�P<�Gp�D�y̻��lVi���]����
~f�t*��j�D������X&�[�}�R5�����#�Nd��R��/+W6��O�ṙ�@��,��	� 3۠|���69-;0k�y2#����=佁۠��0��!;�%2�,�D�L�*	{h��	� ��֠���
��Ҷ�a�9��> �}�ا����Ӳ΍�g3�#m�����
SlY��Z-� ���d�@�B�ް�U���aX[��w�*�ME�b�"���h��>��]B:���^�l�|�֦���}iM灅Q<f�u�5١G�E��mТ�Z̋��/(��.�����\�1�X��qeM�l�g���juIdM�5B|`	R�0t3�b�����K<L䧰��N�W�����M�T�J�z/!=mVr(/��?E{!�1��-q�"zG 8�o�ur�(ɯ�)�~Ȍqj�"z�� o���E���4m�Fh����r� ��_�rC��WSM��m��	�К��)�4���_��	7�@��%w�4U�Z�$by�>�
m��W���֠�W�!fũ�.,�`�Cz��\ljǪuS�N�(ҧ?�q�r�NM;�)c�n�6�0W:~���m���)Yu���>mM-FR��MH���Yz�XM&��+�>x�����5����\�ʆq�Ɯ�QPpW��z�dwe���U	0q�UR|��Q�Jp���E��.W�s?�_��VG{K���`��>sT��R�z�����@���N�ټbgGpnm��ԍ���%�zӰ���1h��a��t�830Ռ����q�3��3�p�Ř���@�"ϭ���&Ǎ*d�ѣ��}M�ȥ��;�Q�������T��'DS�Z.5����x�x5�J%����
��n����wg�,H�ʧv����9o>d��bz��^�ov>�h���/s���r�fs��.�C�BX�f��&��JIJ�P3y���� � }��٨$�S7���5�Y��������G�^^�r�$®�ON�8wa���-�74 �1��>���@��-,�Y���|?*�?�)=&��6i�L�UFm&���y�4�׮�v°�9�� �]�d0ޥbɞ��B�C���}RGn�X���MR��+h��Ru�ڴ������O䣰��ԋ��ңde���-r 8�$���=��b�P�c��o����w.֩$�H=����(K��d�������[����� ����n���
��`J���Y<r�}C� :h��T7[,1~��7��u:�F���hd�V���'k�;TV��@�����7�k��,���mh�p��*)]׋+ܧ81�����n����M�*������j8��~\.U����S�&���l�`����D񈆭:�����w�/^/[�zV|^@3�0��c:^��P�-�!q
' ���&��p���_ P���<<��|��B�X�s��ƶ6{�N7h���V�?�߯;�l��#�Ο��ka��K�r�w�����5�9c�h��>D��a�O���cu��;R�y�3��-vfƢ����[f�y���)�Z��������ơGf`9����7�m���@��`r�9}D
ا��6�����T���6�����⇤!ǑU���y`�*{�ˡ�+(�|�m9���XBm� X��_޵��dge�c��D_��K�s�Hp��	��3�̧�0~Ή�4��ղX%�q18�SZ��i�g�;b��5ȷR�y�e7��{~��J��J��U�aߛ��J�D��q�o����3bY�ao���Gsew.����:,�S��bk�ĭ���S٘gC�˅֖�Ψ�pFx�:��T�YX[�S�	�ђ:��N��2��ݒ��Nֳ{���O/�5]�����G�.ؓi�)$������B��?8F��0��7L��q�^�7������h��p�߲�M!�����Ų�X3ч�8�X_�;.�J�����s�����)�y������t�}Ԅ��Ūǉ6�Jw�����Z�h��*�(�}3na=߫����Կ�E�y@6�M���&,����A"4��1�=o2��B
��}\.�fUb�sE4�&1��@#?֦�a�&���k���`��6�df�6�%� 	U6�
Ej�\r�<8�(�"c��
��SG�GG�x�w�9���Ke7�hHF��+�Pj1i �*E�P�{��:. T��Mz*�D��� ���>)": 	~���=w/AP��
D#�c"�:��_h�R���F�eV�X��l�I��ߏ�'�ԭV�:��.�i���`�ߑ<�:%�$xlf�E/�����:�e38�J;E��J����{��MM�C�X��b@z�P�����������X�����;(�Y:�v��G3t��0�L�$�^�"�kK��~v,�+O��Ȇb��`�`������MC+/1�M�F�IJ/��@�g�ކ�5�AR�Q�Tx���͉]WN莙qF����Tx�]9�W�A��`�>�D�w�ӏ�n�CD��`�:RM�@�.Pb��
�1ⷅ��X�Y�Ȇ7]��bu�J�,��C���Y�7pۃas�N��c�P
F���?h�H�S��G�[�tCe�h[8:շ��H�~Kc�\j]�f���+q*H�!��Q��2�L�:���8Վ�R�����i>%^�
��<�{06!��Tzၤ9h�����·0w'<��'���`~���Q�B^�Lb`R;��:��yda�v6E�����R����M���9���a���Y����S��>0��~���ܛ��G`-�i]�6j���a�*%����1h���	�(O��G9Nd��˃��Tf��g	��c�e�N�>��\�c�k=���P1-@��X}]���
G��Ա��?���l�/���v�+[����6݌�����Ջ��u��,�a(�g���D�%�@�u�7xeRߝ9T�.�	�@��	�h��bŶ`�:u���Sr��*�Rm\l������^x&���K��J�����
�2�Z��f��0��4�ҜΨ������p8%��R)�����H
]f�	2�*A��og2��y�w�3�_���}%hP�x�6��Pn`��f"�^}��Ňƌ���D�U�����,�F%yo)9���M�{�:�k�=&#��Ͳ��&M��ߢv7� �i3=�% �l���Đ>72����W^�ы�EXX4��C+{�z���f�H� ������%}����%0>;n��x�\}��(�~ ,kdK�t���%M7V���W^�n����ehY��\��z��̕.>R,Kg9`fV˄eNH�[�u�_L�TJz���Kg�0�E�&s�@�E8k�Il�%}���A�i�3�Nk�]�7$��Tf�ǽ*�N�%n����Y�s{$��)�ϒ��͐����ʺ��2h�
�ah\Y���,������K��ո�ya26��6�h��R}� ��L���!}���x�x��/ ��I�A�����o<�a�Ѷ?C�=�B���KYmvwe��.`[�\UT�١be\pW��x�g=�Ws*�0o�z���ʫ
���/�����>S���G��1on�X�:�l�kq�*�����t��s���Y�i����=�� P�S,��y����g.����m�jy���/� �O·��q�? *��g�D�Aaw��z$p1х6��@[�m|����;�ť,����B��eܫ��M�c��4@�t\�,TF��_���e�,��Ra!¬Г�v�iW��ۇ�?#�*�q�k��MTU��'0��Y��~��9%?wtDoP=V��K�3\�����ۛ��{�U�a�1�.?�Z���ur7z ���!;�6_+�qGLǗ�D�^��g�QY<b��¦��]7�� ,��%�)A��T�w֍�,����~͗�^g�+rAs'�-e��G������"�x�bg���ز'y�5���(�4���3I�@���!�i�c����!�T`�{ͩ٦�G�_�U�m�'�Q��V����.8GM�X����'����[ K�=h���h���*��&�F�W�N�1V�6�Xd����^�&�X�Q>�t����h!9�H8\�^ذ&כ*�N�yů��4R����[ N.u� ���rX���üBB�75���˺�+�
Ӧ�)��7dmZ̦b$@�XA��ʪ��1H*P������7�M�5Ն\�M.j,t��%�=�[�����d�-��Ewf��;��),6�-������Jр�v�a���*��b�i����H�󱄧��@�����h�E��)q���hb�M;���#�ԟr��E�m�=����$s0i����)+ו�Z�덓�����,ae-ᇉ��e��8Jq��������)�����I���I�:�����~w���3�N<%�h/�ꕸ����b�~�XcXا$Db��ŉc+%T52�B�:Z��Y{Y��C�kNطa���S�6�^�C��5WIY���R���?�OJt�6 <4��6���`�� ��<���C���?Y��� 2$�2#4�	���w��~�����d����e�t�S0V�V�H��}�ߐE���ɤi����Ʌ�=X5�2
�r9:�LqVH�����XN��/��F�ҷ��(�NfOҷ�;�����6߻���%E$K"J�(�;��gq@Vm�^�G×ۼSMx����W ������q��hR���EM3Jv���4�2��5ò�K�d�'`zd���LH�<mpn�)�R���[�I����FЗ
9�xH�ވqgWd�Pe���=�34��1�;;�jF���b���s�}�9����L!M����Y�X��ݥD�6z���T����� >>�U{�n|�N�R��O��o���7�C���u�\�� �P�����A�AC��3߻n��R��n���V�ׅN@�O�l� +Ы'���skt���J7��-�ۡSޡ��;��h��#�)��s�[r���4O�{� _yB
 RF��rG�"S@04�W`��Sb9^'v��T�>�b�V�����@Mz��pJyg��z�6�U�3{�j:��'�п����*q��_8�L��f-२D��W.� .L/2i�6��|��@Ʉ*׮XK~������C^b��s��0w�tJg�L�� ���`��8�kń��LY��Uf�uOG��46������Ѳ�M��Ǹ�&���ْ���+�k�Z���.�(�o8d7k%��-;D�].Ă*)�⺞�p�!��/M��p������W�<��H�O(� �BaS����-�$PS c`�Fl&���8q���Z<�Ub��<> -_�f#x�xz,hDL�d���7S�Eޗ6�Q���)栱7�%d�~��g��c�A�!�DV�
[�����w:��>��F��O�K�ڨ(�k*55p��7�S�9�:�^�匄#vj�ץWƃu��&��A��z��B{��9yR5B��������o�0��eP��nњ�VGD
aKj,����`����ǒ>�F�t+8��-��B�����P@t�������P2L=�Bnu�:�9��
�u�JHR��0���]��	�b��(h- h*�k;������>-VLUdg�=]n���;���F�B����܃��L�se=�t{�ݘ�uw���P���y���Ƭ��%� ��lW҇o�0���>���Kؽc8�"�Ӄ�E}��͜��a����7]��3�"���hzzRd��L���D4�E5���f���6��9\����S^Fe�A�)���{?n����R@��><U���l�����;UPPcGQ�K���; �I_��k�eڡ�h�Vi���~����O�p���̑��|�]�����o�� q���Ⱥ�*��! �}�|���ϊ��B�Aʚ�u���f�L鏰&�b*�G�Ż��@'�'-1����?�`g���ؘjp��V���7hsԫ��@�=븞�ٰycʡ�$F��>u&>�Z��Q�iV��󞫼d� ;�&Ï��= U�h���Cfӭ=`��ګ�mwy7L��Z��&����9�A ��X8ՙ��_�T�}�"�cY�6eC���W=�!�SW)��B��Q:=�a]l#���]�I�d"���˄u-^�P���S�~?���۾����Y!rt uw0��\u��6
OT"�i�l���&K��.J0��t_|�`tc1�xC��!.PQ��G�Yn8��ƍ����{����#	&F�U�
:�ߏ�C�]�K�
��5�����;=D�U �X:rk[w�Q�Y.��t��X��U���Z�cs�L���G��E�5����T^O�g	�'�q��Ia���G����F�u��WȊ�nq�3�W��M��X"���8i�|����v���>��д��4���T{�0�B<�5i�.1 Zi^>_nj=@���3=��L.	q �7������J�ۼ�&?�D8r���ú��P0���u�xuϪ5����"��O��n@t4hUb~�^���.P���#��)�P��>��0,'�֠s�	nm��n��2���`��޼��c�n 1�q����]��{Fܫ� }�adl�3>:�`F�R����h�Uy�	�\*�����sQ茴�Ho�::9�q��d�j���L��RMH44?��;��;Mk�ޯ�w�EN�)l��G\p��x7RVI��֙�s-�5\��\��uxs�?;-�	��n�^ɤ��t�V}����u���8۝��r��\f.�b{�1&�+?|k�&1�}��R�A�����}�d/@��o�0+`���v3�5���*�|�I=�Fr�30 jES��A�ڌQ`:{��´\+���9��k�4b¶���W��}����͞���
�&�*uAN!�RtuQ���>��\�1!����3<@�"�
��9�:����bO���M��f���Ka�X�;,���b��j�F�j2�2�V�"�(I��t�JԪ�}��ۥ�zdT�6|/��s���2�/i&�C}����˥��Գ�6	)[c�(p��"0Ǳ�
*��H�e�@A�K/%�;[�^N���g=����1�$�9������KT �U��� 4�y��3�$ �`#v�bˏ����c�Va�Ğ�<��{�Ilo�8B~��W�N�(#�&�T��������(� A�^�\��hc���3��R]�JP�n�j���+a���M�x��[��!Yk=���Gˈ���;e5���$�2v�g#]����	N��dH�12��X������gJ4����-@���8N\���$�n���"�z�*�Y�L2K .�>�t]�t�na��% �ax*?��Z��X^���HV����|b��ɾ�6��$�X��/���������`�K��3������\�e��h���/@��A���9\u)\K3�a#-��_"F��%_���D����e�{�Tl�de [+fW��:�E.<˘K:i9���	Վd�(g�w��Tt���/΢��Ì�ƴ�[���n%��޶��(2�Eݼ/����0�
w�7�	��gs�`��5BI�\:-�Hb��N��>NzP$	 (�$�I���f��ș�`�E�Tn�k�r;p��VĲ90��>����}��(S@bb2�{������W�M�'nh{S�ߦҒ�te�"�n_K�uc[Q:1��|��P ��w��ny�-Lqg�ֲ��ښj�����)	��I�@��.��l�I26�!���1=�s{q)�"�Y`��0��c9�^��H
�e �}!GB����;L�N|R�i�A/�S�Y�N��eX �IS2�"*q�'�����vr!��	�Ծ����FGܜ��ή���v�X&�����N��q*�HD�,9v�Ҟ�ߦ�A5��ߖ���Y`3�O��k�9�XMN��sƦ��R"�}clb��CsH>��
���J��{���4\M�k7�3+����&<�����W��K�=��d����=�u �#��z��s+�sٴ��	"���dL���	�#��ӛ�����Td����z!�W!�ukq�8�1>1W]J'�eX������o����# Y~Q�d-��et�ϳ:g˺��MY9����$��
@����Q�?9�-+�� I,�}j`��?��Zb ����'T|�������VT��t�h ����rv�W� T+��	�7\u �t-ypG�JU�o�¾}�Ш|�� G�[�"𮵙n�C��=Xl��G�� Q�ȉbp�0{I�Ƚ�H��Ɂ���O�38�:�4@I�7�&�ë�rh�`����#@|KT��՟�ɦ��=�i�#���At�T��,�����bV�č�- %�3��'~i�@x�r�����TV�6����XN^ƘB?�����rb�v94b����X]o���r&񟆰���J���&1��V�s��Xd�oߥ(\��VĠ�`�����ӥ=��Ǿ7�^a��s��M�i:��N ��H��<V���(ͥ�p��5���尠�������h�=�DG;i��g]��J�Aw�_DT1U��i^�Ȍ�MM�,�ۛ?Ȣ!��Ɂ��p����̄�oεip�8����-@r(6OA2�$!5��Ted)���l
��6���y�ì��>�Y!3�KD����!��3=S8�A����(ꡑB���nao�>\�E.,��ܑ�C���/���>��K�h�L�K�M?g�3#�Z-&Ǌ�W�e=����0�?���^Y�Z�Al�1t;q����.��Vb�r\�Cʣ�,/����+��b�Bc���"1j��i����W�
�g^��_�^��J,K�#��<]?a���b2|��v�R~�|����`fO� ����a����F�a�<��@)gs�s �݀jʮ  �l Ï��nޑ�L*]v=���ފ��u+ƣSD�|�s*��_�P&��k3�W�<��YI�ڑ��5x6�>���,����ec�Q�/_f��z�̮�r�x[�����!�]H��XG%8lk0}�ӂ'�Oq��(�H���{�Uw�Mg�,��x����]E-�.{�ű�X~��k���b��.�����������PհC�ۺ�����@Ӕ*U��{��!��%�(���֣�]6)w�&�͊`W�(�4���/�z�_�Xe���:�Mɖթ��R��+�	� ���Ё).����\�
+���(�B4��,��	�Z\����� T�T*�o�Hw��nA�[z����@n3�汲&9����)�w`���:h���Ȯ�X�l�e�G�+{�d�1v�ͬT�y�ǜ�aP�=f~����=dJO.����k�;��6p��76xz���e����j���FG�W���l���}�~�n�Hg�|�e�o���tdѺ�1W�G�v����R�1a�������4jV/JK/P�g��o.���������ˉ�$/Jࢳ���4ᢗ�Q��s�[��:0Y�
�L���������� ���Owk����X�����|�};�imph?�������D:U�b���%����+pԼ���eCg���_�
~h�ﰼS:ަ��~a��P�U�m�8Q�v���e|����d�"�"CD����l�w����oNl�k�1��=���
\~����o�aF�> l�3xbgB_��Rmq �B9�ݘ�6���ɫ�  �����J �gA�?cVS�V�B.	��:��S�2���Z���+J��H�H�bgW��Tk�c�E��E_��.��Շ���L��-� ��)�Eʔ���[<kwS��wA��;�y>)�p�d[���&�L?��j|�by"J�L�B�&��tJp9�~	KU��I�ᣓx�Ẩ����,S"����ͅ��Q'a�#d4��c0������!z�PF��,��B�|���}����FH`QF�҈C[�F���x�$q(���*Oc�ߞ�
cЌ�*E�ϳ��O�K)`���oB)�J�?�'��"ڎ4Pi?9ix����H5�E��4	F�P�x�~�&�?hꖼw�OV�FM�U`\zP#G���j��
?KY{I?Kd�a<�Dpg.�R|&ǐ5�F�n��{h��
�A��;V���MU��]��>>S�tl�c���l��4_�:�U��ܶ�����ɫh����I������iS�<����Ӕ7������b\��͋����/k�T���
t(m�^s����w��jw���om���r#�H.�\�ľ�4��v8���^F��!gR
G�-���u�v6�
�l]c==�������SЍ��|?q)?�}�&�}��QS�9��wL�g�r_�E�:x.�Ua`��rO����-׫X��B�v����|v4�ɧ{�#�"���_^t�� ���'[���
����+<y��7�ѱ∺�����Ѿ̯ɑ�wQ�G���m�c�9$�@/���u�m��*�В�$�J�F�O�w��?��Pz�R�l���^P�ҿ�����*���~�*��H��+�O-��wL=d�a��vn���4F`��y�R;{!��!�k�ſk h���=a�fo��N�z6Fw���&7��q�
k�����&+���Df5r���Y�[��@ �J�x�̻�e�U+^E��Mӽ@�>�3��%m��:y R���v'�4���7K�ߍ��	�L�t�M�l�F�~���`y�$]�;,=)�:��^5�%&�����6��X�r�r�[m���d�/ݫ�wQ���9�5��L��T+� �?��Q��4g�Ӆ��ON�
��>�%�!o�[�	��e�q9潎�śB�I;Yچ��h���$�5��sj�~W��E����0u}A�[�8�fy&Z��A���ph�vp!r��{i�Ha_NY%S�.�l�WU6V9� �<0M@C�!�A;`H�f���DB�'W;�2�ͪ�r�җZ�M�Y"�zsKosY�H�yfL+��s�Q��(�@����"�f�g�h]`��J?��SV��衱i�p�k�j�3�s�˲��tzm(hQ�Y�o��I9�!�˞�ˑꐌb���Q����HG��.�QA̮C	���HP�bT
A����y@��soS����j���-�1���`���!�D+����O�(���!�0�~�y�3��Xܫ��M��Y1"��E����q���3 {.)"h��
��ՙ�J�4��>l"���p�g��1Q�m����cϻw�Y �0DϽ��~V1���<��';�Z��jQ���]m����7J"�J�)��Y�&��#1]�/�lN��˽h^}y��E��_Vc��Zغ(,��)Ίz�/Ӵ3�U�UO=�����Q(Ԥ�c��K�m�t-��09�=	�UH+�մֺ�1��7S8��ۢ�f�b�
?$1`�ZoX�N��C[ʁ�i�e�w��P���ĴP�_���.y��� �?��[Q0PG�E8�_MICA0�F�E�8֞����A+�|�+&�B2���1��$� D���N*)NfDN��x,���l��k����sGo��`9']"�u�#6��ksm�7��m���H��� YE�朮����	Xl [L����hi(�w�����sq�����+��c:+���
x%�0�E "]�<�Ʈ�]T���bWr�㵌G�l��g���J�_���㕌#FN�C�Q�X�wy�XE^�]?(��=�͑|96x����v��`R����Ə�����]m�.o�}8Y�q���1�V�L� )����cPM�����B�e������Cm�F_�8o��3�0>��O#e���3�UtjEfz�!�j��<x5Ik�e/�A��^9�����A�o��*�<*D�M�+({?��Y^��>S P��v�0h6�)ω��v��L���o���k��xO9�����5F6ۿH��,:ǒf��L�f���"�GF5��B�K�6~�t�� sm�±�����v�η|Գ��4U�we�:��2P=���'�y��3y��L�P��,������ɐ �[�	73� ꪝ��ݔF�R��n�h>��%:���Y�9ڕN4�VX�17q�̬ʲ���ҳ�_��4���k:h�4�WN��Vy�Fd�#A�X�ҰF�tOP��ěʆQ�D���B��Z�*MB�1���P����Q�}����3Oo���<�ןOfE)cs�֘�Fޟ���m/Q[�����d�Z��x�)�(�6b�\Z�D=y��@.��g�whi��H���Ib$fL�ְK��$]v9;��l��yȭY��h����ٴ~K�b�;ԅ�U��Nvs�3�h$ҕ��ǈT�H����:_�Z����'DH*��N\FO%U๻�s�
��5�%HϢJx}t����/�1QY!�G=����Q3$8�O|��)$�4@\�Sq�h�iz�9J+E��YC�^= ��[�S��P����L�[��xR��������n���M�X���N	.�W�R�)BV�i˛�� 
���kkA�O����ap��L��}Z�#)��#�ͤ��0����1�IX���|Vͻ��<׮{~+���'��d
�9k���l�o�ǟ%0_q'H�6QI=��Hz���*5�BM,3��m�H���;��W���a3_%�FA6\����|�oQ�K1��>l��>�_K)ρe�R9yz����vf� �I�~���@X��ic�[�:�\L\xr�z�2R>�ȷ���#�Us4+~A����\�/�|���g��$��E��9���U;�&YE۳<�>��J#�vۮ1��$��{�� �#�����G�E&���t���2�*�]%^ ��!Y��
��r���s��v��襤�� ����S6n��(;���,�ܗ��+9��'	��+�K㓴L��q�t��nǯj�,��/1�M�ȗ��ʢn����a{'�P>|/�삖�,H,��)q3�VW��lФ5��AcӛR���ʁ��Ӗ�d�0����%
��F��H���u��÷�=�^.1�X�L��!L��dL�g���&<�T���5��M�	4�\A���v��~������ �E�oE-u�/~zY��b~\�D���4e��F껊:�s�h�����lw2۴��g��Br��۵����˙��]��i�Ԧ��JSYMR���_f$��x$�*:w��#%�r�"�B��FdZ�h+S��հbQ׿�y������_�Lr�U
R{��)����T��L'q�ږe6�J��1YI���y����C���v����͡���W�I��$Ȇ#��N��~Y��c��}�K"3m�3�	����
M�\[�a���IF��� ��ܺ|Oy��pY5�ὼ6����HƤ�zϽz�<��ve�9Շ��Mе��~2���kI
z���ذ?g�~H�	�%�<��6���og���� ���oj�m`&�3��X�|m�xȜs^��e[`� [-��"o.K���B2�[��o�jzMج4}T��k��`��E���2:G��l�<H��r�8`�٪ܺ�������4�{0B��Dnc윴lTx����&3g ��M�+j󨋱���i���sÐN�.�~�B��XX �!�7��n�oYe4����@{�͜���=��T'KW)9e��)<�9�hԴ��H�
���ܘ����
�Ӏ����ौ7Ғ�^�EƄ~\/*�I�"=!���Y����i�ӬPn4�fʂ����yo4;�n�oJ��\��C��)�F(�/����9��xB��z8D5�:UHZvwC9Ֆ�(� ��y��M���d���1g} ��Y��R6�?�U��nf _9�����\�l
ȧ�e'�*�2���*F\��ٜj��d\�4 ��	��T��9�z�Q��M�PG�=i2_��������^�3Կ�W�*�;�Y��0����7Ĳ�0Mk	���.�f�t�zO��k�W$��4J�9����������-f0�XLX�)�i��ˌ۩��*~,��_E,��m�p�O���2�G�1)���&b��-+�42X��4� �Xt�&hЄ�2� Z�Q�%���W�}�匥�K��4�<<�R�;t���� 	�����z��OX�r��珬/��S��D;��>���[���`��cU'��Jf�Ы��J���v���&Q�
��;=HIW�y�c?r$i%9�e�Y��Z��P_g��H�tǅM	ư����<d�f.צ��I�(G����<	[l��0������m��.�����H�Xe M}Ts�%�7�\�A@ŕ��@�_�Z�qG@?�?�^zt�>%I��a�Q�7�F�p��s���2��q !10nz��z��2ՠWk-N\�ӴրG����iw=��s�=o�0�x�S䓆��[D��߭=������$�q%,����/�F���-*���wp� %�߭G|H���r��y�d:���[m5 M6�ѧj���}��>�G��kW�xo�k��-�a{�Y0�_��Mq���jgl
�%�Q��'�ˉ��&�em2��Y4heăLB. �������JM�b��ܝ�}�؜B���g)a� ���Էl�)��s��W�%����L+)�5p��]���!ȸ�/i�A�с�9ן8W~��E����٢�y`��@�l��i�����q./"�I񛁖�E�')������9.�-H�����_����N�f5Ѽ11{C�07�l^�#I����su
߿6�����1J�%�a����$V�����$<i|	�7_����ʛX4�nٍDف�N����_쳻�ʟ�.�z<�*�$�S���9����a&(y�Hw�n&kM���1%��i�ܧɾl{8Us�zw�(��l�=��}%"�����}��^��碋T;��~�f�=�@EN�����T���X<�M�i����+�r���W��iwvjYR�C��`�B�-M)���na';q)��Z]��<��ʦpyk5
�1&k��@a��]��15j��J@���9�̅+�.U�5��@�a(>��lC̷�B��ܞ�;�_[�x໠���g-��OBM8 �`��Z��8.����Y()5Sޓ�>���C~�6��߯jK�l���]�;�rh��t�R?�Z���RMa�*�h���#N��ݗ��p-��i�"'��h/h���ƺZv�< �>�
���YB���t�䈴+��6ډwI��}�\N����gp�h����z� ��L���f��F�h����Lm����?Ԙ�XJ�3zE�e���F������m��HET������Bi[v�}���QH�8�Jg�*,�Q=B>����~=�l�H�M�AY23_�}���Xb�����P;�c)�Z:�2ِ1O"��?�����؆��tD�R������mg�qQ^�߻ȟ��t/,d�|s��l���]�cskda�A��}��.���)��x�̫nL�q�l�i�c��
p-����>����t��O���~]�\�-�RE���;���~ť�Y�1Y�ǃ�RO�ձ�G:{��3I��4&U��B@�t�̇5Ϙ�\%⾡��m`߼����3�1B�%*�#���Y�E�n�\�D�K��E�[r�b�Wl}+Ze���5M!	$ҵ��94�Xmؿ�.�=���P��~BS#E?�d��43�V��m7�%1UŒ����݂X�g��\}SOc��K�>|�q<��9�-�g�����������u^�H_���6�>7����?��QW�l,*#��*]w#��J��t�36C����c'�$i*ޜ�n�C,u�C��d���]����IXɂЄ��qͩ l1����{m@\rm������G��@�A�0�R(_WR���O�<N�lmk|M��u�7[�ƚ��.�V0���� ���N��$G�W��Kؿ{O]Ei%v8��(��p�������4�������(t��xZ�?}nG��_lV����Ϳ�cѠ�EH,�EbL-���a|�]$��	��M���1"��t�ݼ�K8]w�O��#�����$�a@C�.{���@�z*��'�q�]�]E�5:�`�Y�]u�$����Z���%�R�_�_�@�P�U:D��N	_q�rɷ��.���݅�x�*�(�X�!����������t�!�vF�}��b�g) �z
 �g�wg(y���Џ������*^�N���p�M�����qT�����~��4@����/�=���i���c.$DiO�'�� � Zk0h	���_�~7>�¢��]l��{����]%`��J�"ˑ=ȲĘ�q�����1�Neބ�Y�@���."�����y<��j����Z=*������{F�Eԙ}�� �3�I 1�d1u������/=��d
�ք�.�@�^�u�bu+��9W�L�O]��ce�39e��<F����@��?$|�(S��6�S�Y�)j��6p�;gѿ��Y�����X�z�v�*�3�!�{jA�`v�R��l�v<�1�JxH��r���?�c/�3Q��׎A3��!����m�4�:�����1ɒ�X��� ���?�}�P@9G����_� �ݏ>�ů�j�r7��UFf0K�� ר�P/�|�6Cp�׊����X~���M��c�k2�T�R\�Ą�T��E0��oΙ\9E�p;�ڼ����5�nʴC�G7%̸� eEI�R��rL�T/8_ �1-<h���/���g�6$fb�nc$���ѫ�^�o�v�]�c'�b�!���[��؋��D�D7���hg��x�f���4�u&6��Ъ�2�>Jm�Y3@��ì�Y���7[\j\��ɷu�K�P��`k��Y!N7���2�����ٖ��3K:�d��_�I������&�PF��"TEe���6��;�EZ���;�q��*��i�o4��7��n���V����y��k&H����+�H2�;�Yߺ�ݑ=�����f,{���~��ǭ���x
���k�A����r�=�3�B�(�X͇��LoOH5/�@��6d:?�*�.��[��q{��ݏ��|�xf���Qr�Y)-��~�;��<��-Xk�8CZ	���3ħ���R��2�(�3х��qDJ��5��S���M��zD�)2�z[�L!���S���&�UѤ�A�ĸ�ǙŃ��Ԭ��Q��]V��b�J��!6+J g�H�����A�moY}�v��\����ـ�@Ʈ�C���E�l1HY��|���'	�㊨~��+ ���=1�w���baca�bɂ�Ⲅ����S���Ty$d�d�8R$�RAlH�l��~Ϭt��>��*�[�Rj��Hv ҁ���Ŷ��I�c�ڣ �f-�d����'ʁt���g�����,_U�Hط��^#����B��'���3�Age�K�dr��?+�ܬ*� 2�X�L�m�Sas�L�Mh�艴y��+�k�6FJr���=�`n��2�������ia�7�b��'��j�:1�>+����!N|�5zR��]t���ϱdU�T�hY�q�ڡ��U,���S�	F[��-{���1@f�:to��i�u�~9��X�F/��0O��#�a��p�зnso�਺��EBd,���{y>���T���|���;��<���N�EB��Ɗ���&�|��r�|���ƂXib�Ў��䄊�B#�k�gm��#��')�v7I��/(_w0�f��+�gH��u_�Lv�
�"wQ
���dL6P~�;�������]���xt��RRݟ�)�p�B+�g���Z����Eu=W�χg����*wnă�UaX�b�����N"���L�U8��K�R\�z��KK����D�{Ѳ��Yĉ�pF�D�K��/�#�l��;�^7�$�~�3g4��x�1	mQ�^f�Bt�Su��1�C�%{#��������UF\��j���ʁ�	1�N�f������d-����ؙi� �)�T⾂/������3uK9�A�i{-L����5�
���R�����Y.���<�QI�Kų�n���:Q�ثW�>�6���G�΋�����clcR�άP':�gG#��g�H���T����D/��7�&b�(i̐_����/w��|E)(���@ �Z�РJp|���p�8�E���&��M�u��䠥�OA6����9�����Ѱ�A"`�2��l���m<�xZ=�^���wBGh���tX���.ID�_���.�v>��L�<A��D���1�Y6���M�I��G����yUT�J���,��BcX�S����g��)���8�R�40:�i�P������31���C��85/S$��Ps��m�Af/��#�h�V-,οE���}ǵ��lB���%��V/E+�b$n�Q|Fe	pI�P��T]�?v`����F��.�� �0��aF�����KJ��:�1��3���1R�`�h�k�e���U���2�Eد
������}�
gMqO�vv�����x�Dm}���O���E��(
���ޟHH����H7��E������d��ʦN^$����;>�tP�-�>�¸AL V�,��i�}�Ɵ0�By^h�T��|\%a��Ńn�����w�TyN��w���v��ze/���L�֬;�?d~4	s���"4y}�am��z��/���B蚸����;��@T��\�ё����xD��-�?��Dח�c�i���?mĜ�M�aJ-~}F�p�g���oM�p5'���`ZB�"�{�QMv���R�:g�w�)���5O�����8�J?q���}�@�����v���3mZ��\��O1M�*k�ID�"I�������x�n��]B��{eh]�G�R'E0L�DrV,�e��W��Jwa$��x3�6�;\T�����f͝�eU�,�a/J���:��Y�@����*[���9����O6��r8[�MjM!��q��mq*�]���֎RFIt���K��+q|
�}�l�@R��e���U���leF�6sd�ݐ�<F�\�sS(>�%�['5j+��/�`ON�)����uG)����_f��W���7�عʻ셊u���r������#��Lv3�f�~�k�V�[��x�Cʽ�=���1�`V�4$1{h7�*����Mu\P����necv���x
]h���c��i�s>p�,a������v���/���zi԰��6�+�ֶq}��!8 ��:��]�#2)Ɋ�}���������w4ԞK��#��HR�� �J�8�Gw�ڎ��~H*;���VAɌr:N�>1�N��Xx���'vv����g|;��N�ݏ�ޑ*��!��J�������N&ݝ�@x'0��k�?I[Ƣ�&O��lF�@�~H�	R�i��NA|��@��1��&�З���K���*{�ɭ�Z�oi`�v��:�d��bb?�-���8�1��HF>�]�r&�<� �,#�.� �$ģ'@]�,�?{9%�
�Q��%�v:�9R׼�t 5t����Ms�y��u%�p<�ce](��J٨EL���A5���������aS�^�P'gOJ���͔B���[�8~l�3�֏S�l������D(�އ�SH ����"P���*3��v�4����vT�����Xٷ4��4��Y��,���ɻ����ɩ�2�B��Zձ@�gu����'	��D��+�.�H��n�&��{��O���U���4�G�Lsq���O�z}<��Q)��N�����������a�&2���ȴ�_�:��;ڏX��ߟ TW��]՜Ƚ	��G!l�pC"$~i����^�Ux�?�'^��U����4U�T��t�JaiLe�S���ݬ�\r p8�����3��q��2���o�װ�N���#e���qR(YȠ��a���ImF.���V/f�{�g��ݣW`X+4"q�����{")��#h��D���#���$rQBB�<�� ASؑ�v��Ț���Rv1��r�MK���`y"G����˒I�ׅ��d���f�0V��i�G ��;�#<3]Kg�'��o�
U�ŕ��k܀�Md�E������쐤G�.d����i)c���R���hg�z=��S��,�&Rں�Ҫ�]@'�4�nE�(0�;��QfSx=�%࣭g��P��(�,�0���n��7��%�0ڀ�o�I�ΨNvh��b|"9�~��y�|�ֹ�`i�Iz�=���x:i���h��y��X��2?�]~�F�����bv|vS?L;�^�Bb�"3�*�I���y�9��B�Ψ�����ڵR`���k�J���Atg̴� �����J�=;�P���O����$������p���q��_ƫ���@��TA����G��s�Z����F��6Jůq��w'x"&�^/ϛ�"sf)�Սס�+�'_�?�u�G�R;2f7Y�}��5�TMհ����=f�	B�G�N������4�K����b�x�ٓa����tf=�1���X�z���Z4'���g��B`|��`)�/+6U�4�r�;3ZK|n�2 N��Z���S$�eZ�����R�P
Fv����(���S��+R���afi���퀶e���QIn�fT˄a7��i��0Z d˄��%2�g�'��4��&�z����󕃥L �"]��J3�rJ�2^-)�^��v $ﰹ�6A/'�c���1�c�:�Ί6��[�������T
0＆��A��ª����ě�?6U�/��\�O~�H�z�Ư��%=���p�ۧ�b�R� �q����k'�oL2�-��֘��������^Gɟ:fAf�y�&�+�����h륛D!�����nUݎ�C�¬?r|Qs��Fsgl�(���&Bۅ�]���0� �D�� v�:�+�f0b������ZL4����>#/c�2즇ˌY��HP1�f�~S­D|ܡ��8nFqΩr̮�c���C�2f�?x� �xyO]8\=%W�|L��EDkɁ�;)��/e�(i8�O�.G1i��*U���c��u��{pZg������O|�	�em���D�v�|qe��5�=��Y{��~�H�(	}u��D�8�2����Ru�*�$��"�t��g��: 9 ݡQp�;�Ra��܋�5�Tt*��x�h�"�-�?"r#��>��-�����e߰���d�}Y%r�w�G��ʴK��i��y<�����ږv�����N:p��} }��al(�a���ɏ���K:�i*O�ka!O&���i�c	�W��\9@�9c��.1�n�������EfӖ�8ܲ������H�/V��l���,ٗ]Ǒp*HuSj8B�b0����*��`T���6��s���6���ro0����)����,��n.�,+�cpB���E����ǔ��?Ț})s[�yul�o@+ä��%I�?�0���^ܥ�H�}�-uudF�nbOFK�x��w�� 	� �>:+.VmC����E	���ճ������MK0O��:D���T:�7 &���Y����O�n���|����hT��&��ig[����CT��J�����C*����E(`}.��܌��\��?���Iڌ��J�a�)p��"���ˌj~�}d�Q�œ�`��M#՚�ʏɩ�������/�������^ �>��S�/�
����pʛ��n��/�j�7���#�l�ّ&�.ׯ2	�lB��i�}���i����bAF�w�/���0`y+����T�[�[٦A���e�o����ĚA���?{Zz|��Y��ߒ��9���Pe�ͦ
)�[-����z9lg����C��-Kb'�C��Q�_k��V&�(K����q�`���[U't�QZp�+i�I ���E�������� �s&]�d>�l��;��������0�N�����K���z9U��9�TWY�r嚭�4xh\ǗIZ�6k�ͩ�6I��^fH�`=k���+Xʘ��f���e�J��^���u�u]�C�/v�c��,�>��l���oP�#ghu�o��_k�d�<�M�|�w��_A)Ar�f(QQc��4¾���"���#�u��,��J�`&��������X. �!���GD�iDU��	 �#�g9��{h���Յ8�!Ns"��b� ;�������t��D�e���=�k:�����f$=t屙h�,%1���T�|�K��YT��H��%��L�hb�HG�����@{͢lc��L	��|B3%F1� ���+�ZƠVx$��4�>��8�D'���>�ϡ-�Y~��K�g���/�.�مK4X���h"��KC�F��8�S'�O�A���sqUd����M�r�{�]k��Nyb�
��GF���z*:*E����]�׫�$C�c�Wx�W�5��	d}��VL�Q���,7R��������2�/�ݰ�^�	c��h��"�>��Պ\�K���]C�_�ك�ЁZWƍd�gZR,��`��Y��8�,q����
��n�L���\�TA����~�q�![P*�.,O~��GC��q:��n�p�YC�v���q��J��?hy��-�׎cf�..Q��b�x��ۑ��ŭ�T~��FS/~��#��u�#鷹�{t#2�?�Cx+C�N4O�6�����`#2ѐ�@�;>Fw砈G�����N�YF��xl�)��˾� �K�4�z΋O=�&�ە�,�x_ǂ��S�3-[����1P�d^{�RY�.���q�����w�c�@H/�?�ׄc�
�:�;���u�9r���?�aӭ���F~��� nW�=��>�ː#+��ǁ�Dޫ@�+B�\9:��%�d���i�;��7�k����:��pLW1�߮������r�I�Is���̙F�����!Sn���t��L�`�в�l(COjτ�*麋3�X]�;J�jJTx}G_� ���sʠ^?u;��.��5'�~7�żhMT)�fBs��zvPN28�e�Ʌs�rh����$U�^��4HG��n�����J( �,�x\�M��9co��O��󸝾�.��/n�o�a���h��]��_/��d0ՠ����WrH��`���,6�x(ݘi�;��wê��ď��a��流���%Q=�Z�u&A�
�V�ސPw�ݻs��3�fK$1��ҞE���Bɇ}VR�Z쇞��L� s�!�	m��g��3��P:�jZ���S�G�#e���v���C����kǆ7�rq��%�z�v)��� ���J�2^�L�1��ЄJ'��t�;�'��1kٶnWN� �S�����\�J��t� 
��Ï�w~t}p���y��dC�`�����(�!bAUjjBe�(�}��#������Ѐ�_2�:k4�t9�M	+{k�J�¥�������<���!�wG�_b|̖Sp�������~!%U'�9xr�U[ QI�ґ��wgŜi&��Cx���1�rJl��F#�H|�x��9�)��?D�$�}�8����}]$��!�����.{Q),J������i����bǕT,����,�7?�����[�ƽs�W�n��*���Vc}U4�i?MO)Ƈh�&8���<���ĩp�j��ĉA+�_���\:��e;�g�(�N8}upF{��G�ӯ�h����|�Y���Mln�e
�m���F���M��w�N�����-�X��Բ��H��`'�7����L&;̺��덊%��C*���@Yd�w*��ܶ>()�\!M��f�ZoB�(�;SB�%D،������_J��bְo��S4&j�H����9�!�A�a��\��C�*߁NS�5�� �?�_}�l�0>oᡇ�B���_�� .�������1=G���JfDֈ���h$<A�R�d���AX����Y��ߤa��"�AO�c\���:��ů��I��J��݁��ҙC�`��+O�O,璴 Q�r˚1��s�K���U:�i��[� E
�P��T�s���Tr\�t5�d�D�}�H�j�u�5�/�F�РA��p1��-�0�K�Ql�	���v���í�Q����Ҹ�c����Лgb�hN۽�U�i�K�X[*�2��!�z6�2�F2�0OG�P��f8f0=�Z���+��O�0����?b2��F�+֐9:7���	Ã���6 �6AȦ�j�0���z���v��	}���Ul'褛���ੲr�C�~=h���]�U���%G�s�%b�L2�uY'd����{�M�%,<�0����9��3�w0�nU��7����M�(.\c�/ЌEfpKAp���6,:�oM<ޒ�,}.J��`\�"��v�&
����6��ojn��� �'��QZЗ�I?Y��됶�t vfZ"Ԧe9ʗ���}ܴ���$#���G��=	�`aBv~�D�=x�]F�;�l0�'*�k�"j�֨�
���%/Y֕`eM�� ���U릮	�H�?F��]�!���#f7{�&mWN��-X��1����~̗a�cC�,��:���3������t#	sR�qe�K��_�\r;������L�3�6�%u�~�$𱯲�G�ߜ�|�;{�u���d� ��p�f��>&G������^�����Ҩ�4����\�\f�j��#�I���d�,�>���2��$�1N�� �g�#�9�J���W�N޹�вf����D�<�f���'�����#bV:Ő��"5��R&�`�WbzB��1*��"�� !���z�x���_W/������Œ�����X�֫��[�˙���@��X��+g�z��I�^�!��z���Mrf�0Ɲc�t�P�U/�||%m�KګB��tA*�zI�)c~KFaԾe���5�/�0K��}MWT*Z�LUA("�"#�޶��'Af�ǈ}��x��J�IE���q�9(?���&I6�_�J�������pp��@j�j:��t*dL��f�����J�l��j n�L׼/6��ςIp���A$Q�PY�ćMOv�]���8�>�x2�';�s��"���q��R�9U���ڃ=���Ν�0�	!ѐ����Q�������5U���[����T����%��$��,D��I8��WS���N
��pK�q�Py�I0������$NKO���<+������^� Åy �*�qb���Y~dL�f5�<\2�4�*����夔�vŕ��'i�:��!3Ϗ�Ԃ�F��j�%V�a���d��?a�V Ƙ ��}��/���a
�V�P����]|���|D!�cW4^`µi�k�����奞}��g�2�Z�I6y�n#���8@׊2�3)�S���~�zhQ�AH��S���HMw9��ɗm�b�ʙ�e��7we����cS?c|+n�����C�| �?�V�R�T'�2"��rNØ%M+���)F��(�N2P��� ���nQ9�8�e>z��<�7���o�}������nA��B@D]���a�F�`y�}1�K1,�gQR�EdN/����2�gI��ƻ-J�΢F(�����
� Gh���W5Fv˗�Y�uO�|q��k��E�G���̰�p&��(�&��^��%��������>;�B	�_��\� �W��3�դ�� �v��­��܂�b{�/[�����B���9���Ҽ���o�3#iaKj��<yɣ,��a]Û@�xU��>��]����>)�)��Dܧ����҉�x��r���P�� @���l��O=�HɃ�/(�I��x9旁C�������O�.��m��M@�{�B��U"���������Y�`~E�͇!w|T?�Ng���>,E"�:	a*�����<ˢUYەj�� &!v�QK���*0��ʶ�繀6�%�����sAU�{;����E����$B'(��UX�K�Y/[��>!~>�>62��c%?�K;����r�uBL�����[�������x[ �|�ץ�kϕs�Q$�a�;ޚA��������o�����Z���+;zA�v�U�`}��?�E�
ǥ,)}J-��",�B����WgD0|Q���*>��e��\���t��;l�b������=-e=F`&���5�L�|3�W�Ty 5BPn���` 4�w�,�Z��	��*	b�y��ñ��f ��� M�!��1��T��#_-ۋ����^�� �J	�7�ǁy/0�"<"��i�AF9��������5���X�S��k�S7�'��+*�d|O����s�����>[0cB�q�;#��^J{V�.!8ݤÿ<�
�o�>�h���8��+�e�"���W`SP	Y�K�F1㿫���\�}Jb�7�	���uN��-�.
m��H|]�8�tF^�F�A��2Ȃ�P⺪��MU��N�/3���%�t� ԥ"��P�}pkеpt�
~��	��T���̇m0+��Vz�Ny=��C�y�U�iF�UP�ߩ�������o���"W���f̀����]��=4?Bn+�M0�d-1U�@�&:s�ۚF{�<(��:��5b�>�}޸u���a����`�����3���[
_0Q���k�p~�NW��mg�V�r��E��bU��d@�*V�y�Ί鑧0�۔�/�D�q�B�\G-F�Y*�0n*T�Kx�yzw�a4�-Y��v�����`����=R$4_v����:��6v	�'��M��f�5��Yŋ��'#�h�@�z�B�W�{f7���N��k��M66�g!�:�:���ysP?]�g@YG]�dCg���eB�%���L��yjTMp�_�����$�ܙu��ၰȡ�k]��B[�6�M%��vҞ'�7v�Ȭ9�α��X��F��=�N%��S��;���٩��#�f�W�P�1��AA�k�g�8�'?�@s� �ugz\$��\���:�R |�ݲ��dH8�q�	���j�U)B8�>�>I=$���E/c�]����w�/3�{�����(�?^�ȧm�c��{��*T�4�^4�O�'o�udJs��=��9؞��ށSzV�a6^����q[����t�M�^⮵����|n��)�2{�o4���t��I����b�S�6�y����~��3����w��e �}r�;eb'�_2a�Js�0�&����e1m�t�s��L�t��Xt�hū��6�;ɱ������i�%�ހ�N�5��Y���F�_o������
���j�9��|�d�	�)'FY��)ϟ�������N���i���ã@%�vUƆJ;�m��W�9������\\���Q��pu�d��͵;�;F��c��%4-s�a��騷,�@`фt��e�k��F�Wv�[x��u�:�s}�	��D1��q�{�d����,H��|ڮ�~Cn��=��|�T;,�t�V{v[O�(>3	�诵�3)�b'o�J�p��i���`�}�I4�����&�((����e$<R�Lx�*
�v��`i�Vf�ĺ��-�#��vI+>��& ����7�|B����5>��S>�;�G:��ܜ��4�;P��?U�`����hFJ��i(�W�n�1����6�_�3	Ȁ�=\�GI�0�y�Wv���6Ʈk�Yq�3�2�u����s�L�đ�1�_~��vW5�9��a��d��ݟ�b�N�����y���t� g�)Im#�T���� �C���9��v��:��*]�q��d�,�'I��$�|�Ɵ���a��VV�q�C'6�`��[{�[̓�Ĉo"��������
�G�3d��tI���K�J��lv���y߄\R���3��ʾA�����c���r$5(�F�ԁ�J�|]`��L�>�i�S�q^��<	`j#�����t؎][��e���'��d ��~�4I�+N�o��
�����؂<~�~k�N��{
�D-��SL�{���]�5' W��3I'���=��SI���G[#&M��;$��pR���,�Xv����4s��\=�;%�(�Q��N����p�	�E=$�QJH��>p��h�~�x�aM���WUzr�G��J�nGB@��h���uȩ*3<eAG��R���	B��A�a$[D�̣�LҋQN����`Y���ρz�u�x׻��Q�d��� _0vc~
n������zG�����5��A����y5��:�k��6'���ʃ�O �PC�����n��Ƅb���|�?��^��(��0���m1,N���ckL:�7;�����o�hȗ�9�#�:T��k�z>_���{��2�sM"�_dՏu-��L:�����ݻQb����./�>adG7�U#X�L��m��#G��k�t�I$ީM���������m$]�d���ҋ3�2��OW8�4�1�	��n�w� �����FQ �h�4-����ٯW�Ү%�o�ϟ�3F	a%��Dz�h��}$I2BD\Bj�$�C���
�G_�2_��\! 7p��k�!P���~�T6n҃�qѩ��4�pߎ�7�B�e�h��.x��]���i�vU�����#���i_���`���J���z)�-R�M���<��WjB�OQ��6��b�@.($��;Ъ\į�xΰ5�����*�7�
iy����L6��q�ޒ��#+bx��@lv@��,aeC��:ˏ�����U�1Å�X
}�VȽC���[sv�1d��	AA�X䒱�N�Uf^{�8��{�a昰j����[^H˄��e�ܕ�ϝŗ����s��8|;ݵ�����?%���j�o�'~\E��)�§`?�s�e���m�ן���w�����U�����T~�V4�5��u {Nu��{�v(�ގ�nh��=MU䇔&�ڻOE��ү+��sa��?��|G����Xb�&j�������������2����O}=h0�<��2�����q6�29|#$;1�ZQ�9?O�I���	�V���	~t��\��I�S�h?
I&�^EWt�6��j=AF����&_Vi��l���k{�S~ᚌV��XM�e1��L�˪�ͷ�5��x�מ��z�UQI�s.2!ڐ��c]�{�7�CcKE��d�7�a�A�w/�<��/:*�q���e*�w�W�X���c3tE|/xm4�nJnuH9�Joc��K\��`f�#���_��s�����쌄��{[�.hZ@T
�A�S�K�]8��������������;M^��"&%wJ���En~�e�evwb"#�GHE ���{5���M��f{W�����cE�־���n� ta�P.FS�5.�����#�b(�Zn�鍏�i�P�ցc�r��e/�zZ3�;�����c�~k�ήp�7\!�3�*<���jq~�)5��v�%3F�����A���!��[yL,w�~d<4��DRZ�׽�nݡ���9��-��M��c=U=�U��?�ziћ�E����~�8����
�ܖƏ)$����4����t:��[�23+5���7AycQ7��8z����	] �ֵ�쩌� �m7Ӧ6H�YO��~m�����f�9&>�^kC��7K���߂��a���r�����J�������bL�.�焭�������iZ��Ket_#ۛ/u�dJ�e_�������$>G,�3�7Z0B�J��^V'�2`)Օ�]:�Ƿ�<�z�_.��i��C�5��7��jjVt��
�0z�\� �6@J�Ǧӡ]vl�l�����y�V��8�x���J$���{?����L�����U���џ�*3��+�}f ����*U��ɿm� >��*7� \z)G�b���`e��K�]�Մ��@T�hi�f�xE����z�3�~�e!�/� �},:�ׇ�nV�y����Z�ҋ�C��P|qj���JUv��g��؊K%Ă`�'��H�'ً�Ż��ğ�f;��kea%�<�~�ƅ
|�2CV�E���O�D�	����~
V,6�j���D�뢏� �prgA�e%��W��F������]�BK��)��nU�i��8X���Pᯤ���ן���\KV��zSu��uؑD?�>�`�iQch*����P�Ń��2]?�º��\�Z'�y�}�D����]�ezˡ���<n%��K�����~�������@�-��.�8�P�Z�;� �%u�8яH�Կ$����$�� �!X��s�t����-zz$�+S�.rֱ��4:�Z�~�)d��O ��y��=9Ҹ41xkmV���=6�\�CIp��q�@�uMŽ.qO��T�?���'������4Ǝ񴰄��xq�Fh>�?h|_�A�CG��`nde@��Ǧ��O	����q�"Ύ�J}���|5�r�U�A� 	Q��$b�T����}= �R�E"V^o�$?�M���M\�&�I��ӃK ����H1:B<czz9�@�hW���I��8@o�!�>|®+O���}5�,�PW#��h���3����6�����I�p�Lpd�Q�T�2�`'���T�@9g�8��i����-Y^.���oiL�H���Q8<Z8��$�*cbs���j͒E ��=�����qk$iC?���4�JǱ\]yZ��
���O(���{����u��
���B�ޓֲt�m1a_�/* ���a!���S��J������?������.�g9�}�cX�on���ʬ�!c��Loև���v���@1p�e�NYat,�a*O2K�ge���`I!+����ɔ�ݍ�C%�"�4I�=��EVnū֚�l�&%գ���+�;>| ��	��|��)"�� ܼ �˪��/y���t�u*�.���R�tk�JR|s�`YΫ��(*��Mg*
G�;�e����92���������n�M��}_�5G�{�G�M�� �E'����nڒ��z���=�eY�9?�<Z�:o�a�����kl�BQ��!V��j��J���2�l�?���/�C���'=�wp��a2�-	�F�,�ɦ@Wvs���Q7�G��]0x �`VEZ�jm�;�|'5�6�6�B&�R�Sc<t��[ƶ��T2�7è��>n�VB�,bn���5���e&����T��ɚ�t4�H/��� �	k�q����v�	z/��^��;\����ZF L��'�d�YD����Bv�Qc�{��u|���\�8N�APe���-!���
�`VMl��~�u�����-���\/�/u���8"�|��Q���%���Ɋ���=o.4�Ҁ+}��m�����I�ꐅp.tc/߷���bE�xn��)��a�8���O�ֻ'�䌦��1yWu�χ��^9�k�aǡ�����t|5+�r;�t	���b,^�}�t�����D!�0n�u� ��E��T ��C����[��䨩C!�2��@��;i�r��D�'cqr=�H^+���GF4;����t�4��Lt�$u��Ĳ���Xl�Ep�Ld�V.���)��8Q;Y:���aq����n(I�8TJ�g�v��Â<!��&�^*j� ��A��2�}��Jp��hk?�_��A��3�A�\�[##�#� ���|�������Y�ޠ���c>N�Y�R++r�G��&
\��(3�I��":^[,����Y��Ճ�os�F�]Q%��ą�|�N<�6
�È�F�aÊ��@�P�#�Jh�yB�&E�J��Jc���f�2�n���۽@�L�[h�����q��7.~�)����c���_��h�TT�;��$�h�B�vKZ��yު��=��� ��ԕ���қF`|4Ctq?��1���>�y{Nݿ~�׹���S�
�+�={�.N�n����hYʵj�'���c����h��
����yk�ׄ�#���:��4ʩ#�=� �	�����^��� I�Qp�)��[���PJ`}���.??g��V����%�]�K.kXt=�̺�!߁!���>V�l���c@��0�YN~N߻u�y���z��}�z�wA1$�+[:�bsG���y�DĘ�S�ojC�r2��ګ�������ATl�U��p	���x��}�x�m�7v��|i�p�i�e���v��� �1u�l,��p��F�CT�ҧ1�h��F⹕��<�n2�juz���Ӏ.�9�M�c�
�O������y�%m�'���`������9_.-�h����)�P��������V	g�+���E�����c9�`=a/'�ϖ��2D�|��v��/=�5�*9\AV���D/B&��u��"s��QHﲮ�dT���/UBc��\�X����_�E�=���œ�3P[y(�}�KUݥ��ID�Č��[� 7��cWz�҉�ѤE^w}�n�w���[�;_�&'�7E���"k��<�V�����m��v�lǙ� ��#�Vf[oKW�'fj����baV�b���^�W����Y	?|^��^���:�u�������?��
�y�U�i�e��8�*{n��tI~�B?�V�x�X�k�F���핶�	t�$OiO�I&��z�Ÿy�ِO�*�Ro�ϙ�� -�³���I��)�(`Ļ���י��.H���e�nn)�j���~h*��C��*���]L�ͤ����wz�^��J�9�Iύe��V�vl�WE����XR}vY�R ��L8�c-E�͂���m�P:�/m@�I��:�&��y�yĵҊ����1)zVz)n��3�c��f'q���.�c�����"ί",�.��z�>U=������2�;����ӧ?�X��yP��h�Ò-��!$�Vf`EB�-��,!iG��dC>�&��J�ǾCs����H�E�6��}�J�p��9�ϖ"��y<�i�`�{ �
�Iu�Q�+���(l���1ۼ��ɻ�K��]4��C�r�﻽��%y+�骚�H�W��f�q�'~�5R
����"ϣ��D^�������$�.0]�MvyF��l���"���aLo�N�cUk�}�SjO7��`��\����n8E�b:���tD�]�&�O<���W>VlFU�'��-�Uq��c��ϊ	��%� ���@���_���#�]�^��9Z�B��#spj@��̚ �m��`��u'mI��	�7��2Y��$5��p�g�Y(;J$�c��C��t<*��`��	T������ƴ笼�ս9mw: XK[nS�P���P#%�;F^�� �sM�.�<V���-YkEߢ��Z�Z�[N�R1����v�EG�=��>Pf1�v�2�Q{₩R`�X��" 
��)��Ģn�(T V�+ ��qJ\D�ė�����
5�A���Q[F����֢c��	��\%�z݃_�!u_*�d�j"pɹe@��ô�<�GQR�|�Oh#b�\�4<6P�=�W�_��!�Q�^�����`���!+�O��
Hɉ�e�J�Ye�b�{a� ����� `�m�h\������rP��)��>��{ٳ9Β������K��T*	;K�N��Ԩ�l��|�Y���0�m�* &��bD��bjH� )�{!��t'&��7j����.�V��2d&�I�+~��
օ���!	Ĕ�c^����U%�[��$��D��V�{X�@HK����c�S	���!-K�g_�|�����|�u���ٽ}��+8���7}�l�Z���;�>V,܈jq��5�dSs�扵Nv�kn��m���@U|�0dz��I�=�H��([�(��Fw���4D���ؚ�n!ƿ߆.�,�kJӳ�d���P��8���Y��\����S�Y|p�?��,����zm�����*,�9��rI�[ף"X8�`�C��"�jx&� 8Q��k$��&�	�0m���<Eo�Mc����h;l�U{�&#t�x'sg�n��AQ�
�؍�;Ɛ�I�t���]�I�[���m�#&5B4^��vU2��R��%A:z$�~��9�_�jU��lk���~x�G����\���2Fׄտ�٨����IB�.)2"�+Oup48�����[���1qa�ƞX}��t��l�>C˾�O|�C�|��r�ąM:$�'��L!�'��v�u@Q:��l����!͒=�)ֈ�b������L��/�4�L�\����~��2�H��ۑ
OqǨ\q���&��W��K�eu�2�n�2z��r��|xP��ͪ2���M���(��9���O�H�<:2��)�r��j~I������֝�&�K�=P��m��(��/B������]�i|	�`��c�V)(�· o	�8����M��*�o}���n�tT ��p5��ǚv�����}�s�6r�����@�:t�Q�D������܀�pJ7�rٟ�ZBǴ K�K�<�;OQp�|�W��U��:�=��C�2�����5�VKSu�c8åZ;5�����%?�2��cK75�VݠP�=��NI�T_q����֓�F��� �ێ	mXN]�Ϻ�������g&I?YP����$~<-�U����v�ꉍ���FM����ży��K@eL�¥"�p���%�����1���9�"4�e�~O� �o�1�I{V�� ��R5�@������S���x��wR��v��A�5��Rۼ	����}O��H�0��e�R�ː���y|O-���B� �I�=/U1�Uu�(����IQ�Q`���;\Tv���?�(�T��+�B�X�,�g �i�0u��R���|�V� �?$�܁���E�bG�Yѿ���~�?-~.��u�īVK�WN�#�a�E����Ц�M�u ��ה��C	�I9�~U�"��h�˩������e;��V�c��U��?�-W�:����m�QP �.;n����~���f���Ν-�3Q"/��|A7m+��+����.�3 ��->ܠ��]�0��D\��q��R
ƞ]9�Lx��kp�Z�-~����I��!A !��B%6�5՛紺*Q�`6�^ľ7ӱ�,�+HaW�
1���ɶ���t�V��Or�O��{�N©}V�(���Ď����j���^�t;�P���ra�7��U�����(+S���6)m=G`E8��txW�d���+�Q^������B�W��8���:^;���(�[��|��y��^/������wc��߫����3�2x����i%ф�������Q���*����	W��W
��0��~�-�&[��z��Ӯ��/��fX����C�;e�g�6���t��1V�w��\��T��l��p����56�˟���P���-�SR�U��;�e��1�iW�~1���wJq*���F�B�����h�Q�umR~�܄���9�O�l}�Q��������@E�Չկ���37�p�Xs�V9� �!��{���в'5�al���(i������D��p�3t��i�-Qq��n�σ���Oי=`5�9[U�ٟ�<���G���Y���/���ʅ���~l��й4������%��@Sg����W�Ȇ�!� .�ˡ�K灸#r�#�kRUh%TSe���ﺴ�0�H��2���<t�no�}�;H�a���_�Qt0*�E���؝^~F�'�5����}3�C�C����n�}�f����Uw�.7I�����ru%���0	zf�"�̺�7K�M���E萔���b;�/_�/x�����;::�9�Rr�l���4�� p/�JZ[r�~+m^��6�_V��q��l�I�U�E�]1U���G�h>��w}���hT��.%��;�q��?Ȣ���17c��PJQ��F��Y�j��#�V_�P�t��ycE�ڞ��б�s��y�%�hs��l��5]QA\��*�̢�>�k�eq��*Z(�C���x�F�m���W��5��\)�MO<�
��V���G�6x�S�����U$����0+X�C�O�&S�C��'�I�z<�R���E�(�2����7ç���
����`꯼Ƙ��V�uW�l �2�$���2���?+��=&�4���4i����>�����>0�~N���'(IY2$�r����|��b��vZ/��O�Ŵ�T��A~OD�єW�|ҥ(XY�1j\�)i�uyÁ�[�i�f�UPr��%�^�?���C���''��Jbn�����ų�p�Ǻ� ��#z:�x��sa#���_Q�u�k�m�Z�k�E8��H$�5�R��̔?����#ʽ��p|yJ�npI�x��� �8��ڵ��-9�Ahh�ϝ�';��*p�߇
���D�%@��`TB"�zKAZ#l]19��Z��uĤ�����^)�k�М���Cn+[�zJ�`3'�4�����a
ш9�Φ��g��p��Yٞ'�r*μpD��ܛϏ�{貧��ju���?��⏔]�9��L�/]U.���d<���t�(���lhL%@��P�M+F0cl;��?kv���3�����U�ֻ�ޠ�G�D<g��.��_\�C���r�Egx.���B��.�H͵��c�"��<�%�3�8~��Lu�(�i����2�%�����'?جI-���]�o����[P�z���5���(���p���Q��	�c5"��F*�g���5�F��
�t{ܵ����e��Fŀ�V�FS�b�`@Q��l��@�d�����e9c |����MG~�H$�`����PI��i)�P�.y�%�/`�w��-s�r�|��t�љ`!ƙ����>O,�'.�ճR$E�\�J�|�.cF���	��.�/$�!_D��r�D�%b��!������65d5�DR��O7�� Uw�L����N�,n�]�w�=�|�_�O�`���V)<��4b�K��nK��`������}�`������U�a�ˁ/O�Cg,B~��g�\�@��+˕ݼ����xTB�DB�����rց�GA\�/����SIF���A�l�#6&#ў2�j��ZM��ph�yj��P�j������R�8���r���J���5�7����=��$z��7���9pX���S��q�(m�tX��]����5�	���� �a��`��Q�2ań���9r��9��� s������1��q��W�J=S�2İ�10�T-+���U~I+.lIV����1*�"Wk��*���o�Z�a�1���W�m�+�?�Fn_�ѶVê5Y�`��-Ex;!�(z��4�Z$����l3O�ϥE;*�y|�7�߻Y�#�O���0�Ȑ�B�@�C�����7F��P9�'/���`f���z�H7L�v9����\f�<���/C��X�#8�Y��[�b0��w�\�PشŚ�h��X�*��C�T� �i�E�; ��$��.��s�����������	�,n/a@W!�ك�~�G�[� $�n��Rdde�q�bU�Р�¤��a"j8��Ɖ7[ej������-b�9�ψכJ�販���$x)F�	�j��nY��,.(>���sf�)<q>+^.�"�>ױ@v�5	FoR�A}�ې�S���w���,�������l����Gh�~��"���q��|b{�M�P��4������4��Y���+��R��b�}H����xf�TSA�^��r�����,� �J��N��/�f9�SEu�ɵ��Z~�����!�͌19D��'ᆅ�7��qe����r���ˇ�8P���8I�Y���,L6,J+��6b��s�����$���]؛|��� ��<�3�n�V^��Ɨw��j�7u>�"�f���/���4�t&�%ۗ�#_M��������t�����(x�{���'�BL]W\��0���*��5Q:�ȿ�߃�!�9˄l�]�eD�4�ɿ���1��!���`CE��\ޣ��[b�ʶ���%%����Ys�7 o��m�	#��,5B?��5��� ����I#�W��0� n79�gb��m���u7��&6�6`�	9Z^�pRԂ):�Rۆe�j~	�g�+1D��3�;��������1�pX�'��Syn�_B6wVk�Y>��Ǐ��1�nZ�T6�62q�3�Mf���fx^��S��r�I�/�$>����F�F��Ԣ	��`'r�B4|2:��6�����Z1K��$[1I�"���X|K"G���ūf��+�/d�Q���L&���|?S;��T���
���y��p�x�~�����vP��1#>gU5�C��N�:2ʧ���W_�De�}f�ધY�bl/�"e��|�����ˮJ 8�G*���ų۱�H��jN�s�N�N*�|+�]�U��N������&~��qD>߄����R,�˦Ų���������r�H�2���#3���xS�9��'����(��J�������5�S���cښ�qwL�Q�Ӹ@r�����S�I/�8%�W�H�Y�+F�+�/�e�q���!Hi���M5p˓�rb�d*L��@[`,��pR��CYR;K�}�*�&�;��֜�˚wlC��8�d����c���?�d_Kc2s�2'޻~�.���]�ܕ��;�R}��	�����^;t&uhɢ�$����˂���䳙T�A9z~GUx�����M�(�����+}�N5x8�#mSC����
���kb(���K?-Iz�+X۱�nu��q���C*���L������:��M�`���u��*lM�ɩ2��񥢉���P����J�+߾Íװ��(�� "�-������]Vָz0U	[@��"����Y�-9�6|Xlڥ;�zԿ7�����{�է��Y8�xt�ɈL��в;1��'��B����!��0�ǕUMԶ���j!��~_�6�����K�v.�͂\(�j�0�Į@�j�o�w|����R�����z�iUQ�o����_�G�nF0���Xg�����jWioyl�����M�ρR#r+�j(`Iu0!������Y�CI̾��i���z��!>.J�'x&�6�5^��%�Z}w�����W8_o 4og��\�dx���o�qv`���տ�.I���7�.�g�Y��y�H�Cm�"�݋��-#�r8-7S������o�B!l�<t��3_����k4�PkkΎ�	D��,� %1��>g�¨:\�/��c������^r�.N3��/T�&.^�&�P{���>^�}Q���Q�;)q�u�^���XaZe�6@욑�20k�M�%�.Sc��i�F]am��m津>��W����0��ڱ�%:��:��S�Am�hr���\�V��������Q>T�AJRR�Y��]>a,� �7XMm��!+�r{�VB��(�����b�}o�܌���6Z�:+	Q��j�C��$e��Ϲ.�I�}�Br�/�@�^���n,��x�7�2=n_�u����^�L�ܒ�+n3x���i_��|�qЮ��`�v܏7W��ei~�,��O�3>WE􈫰Ҕ�$ɖĸB��	7��t��C�F������b�Jhf~as����Y����W�J2&����V�����Q��xlR���e`�)�bwԵ�)ъ��:ߘ��k�&��m����]$Ζ�+��RZ41��;�ô��U�7���c]�z�B z
��[��2��d47��)���)ǾNF`C�j�����2>Q�͘��ӻ&����	X��*3SX���~J( Z+�y<�e����i�2��y��a��r��T7�r66�vHt1!�śE��'М&U<U�/�R���j�v�"�S��I����ԗ�c�`31���@��i9�%��1�U�F���-2ޓ�j�b�	c]a��{��yk�H��|I?-~rQ(�k��=�iui�ī�6��G(U�1�Vn4�"G�r�������ƺ=m��E�gG�Ac&:^K'�����j��n�4>�GF�6=/=G!;:����o�ZsϫU�X:^��A{U�M^� �b
�j�N�<�t�)��*�dj�E���/!�εJ�g�[��ꪃ�py�����xs���T+���뮈��_R(?ʝ��6���^��wVx��|��Ч!��g:�BG���lir;�B@{`ظP��k����B���<]��1	z��jV�*x7���A�i8M��A?l��Q_~��\J	�v4@����
kK�H�y�'��gH��#r�ځ����o;��>�9�ՇDg
L�p��C���� d����8��e�f���.��Y��� \B���bf���,#�D�ư��ܴ��]��Eu����Fu�)�1m\%��^��h#�o��B�B�Kq���;��Z������-����FZ�-�wh=��T�Rύ�q������O�h�+#�P�f�V<<)q�>����c����}҃=����M\� )����7�g���k!f��꫚�c�3���M\��s(agE��N�)�w}��O7 ��ot*jb\�����Os�gE�*�됡IԶb�;�.����f��^�}T7(��@����0p�O*q��2����ë&ؐ���_�.������v���ݻ�8�Ef�n������i�\ٳ�X$����"#������n=9��O_x��B��X�m��>_�t�_���FqF ���u�?S�Gۯ
q~��E1��e�2��^r-kF��g��Sz�x�%qn�-3�o<\w�ػg2 �|�E�?Y��=�+WH�\s�2(��+���y��a��?���)�)p��k�.�|1yuxf�MO��/��3�E���풸�<�U�Ǿ���K�feq���î�'���a�����i�V~�Yl��,2[�s�=�Z�.���B�<��s�oP����тbrY��c�{u�－5�G��M���Z��[.��2g��ån��ئ�c��$mۊ��jC�ǃ=�ovQ�'���#	�J<~��F�Ƅ䏭 zk/����Ah`[����Wʔ
�Ze!0j;���O8�>_���c�mo%�Zp0�uq&�=���b.v��7��'?�|���};���~�<GoPܦ�έ>�?�.���3��߿��^�P�����Q���A�R������@\��At�b�]g��9��~�����<`��β���t��!�/�m�I!+K��/��.��T�d9`��3��^^�4j UK��[����}���O?��p���>M:8�<{�qFWֈ�@[�_��.�@�M�����e���"$J3��.�GR�o��?>׋���م�8�g��f��7Tm���o���L���Q�)���E/9��%�O����d�C�*�c�����d�[N]=T7����%�p�q�?x���4���D�2FeE�#��"kOI���89W}Ɏ�yd)Vt7��9���~����14�b�;�'�}�󦴂�Y�6�j��*�v��-�������7bg�~���b?%l���c�7�:��Oe	�🸀  ���w3Eӵ�\`��4[�K�����<>>��A��C�Tω̮+!j֗HR����JN�u�}���6�\]_�
��V>��G��+P&m�/�ĚKTj�K��s�u�rY�������p3�&�6$*dtB�e`�s���U�x#��Uj�s��vY��Ⅲ�������;�}�N�W��M'��6���v��i⟝C�B�M�6���%2(���R��ZR���N�!r`OJ��?��-��ly�Cha�&�N˶�}��1���	<z죞��3�-�j�2����'sFsǁ�}F6�#��S��WF\g���'�WM����e�M�_0���
�>�Ҽ]�v2D�?�S�Б.S�PL݆��ZT�sʶ�.�.�lj�Ǔ���A[��9��G�vA`�����ScI�'�1��E{m�����(	/,z6�-��|�c,��e�L{��mps;AB�7w�%0l*�:ͤ��;�#ci�FX{��|颁��2�.s������4�c$��hfSO��L�V��U�.B�D<.� �G	����w�^G��"��"7�7wZ-�Q��"sZ��]2F4��Q���&R�ñ���"N�"���ǱV�[f�.�hRA�K��?�!�N�~%C�2�UGf�V=r�<Mm�#~F7��قX���0��׹�� ~Q�H�n�
':���x2Џ��;_�ɓ��ȥ���H�H_Y�پ�Kc����aK9@d�W�*�-�1�'~}|nN��[Ğ�����Z��ϸ��w��i��T� �Ɵ㱢�yT���9S!��ʀu�14�CnCo�e(Bm;YBw�8�W���u#�U��L��=�Bjr,�[+�����c
�*��B�(j'燿�r+����1�_����u�����2=�gq�5��@��`�n]\�w���P�>�m��f	P�l������� ́��E�w{���oO�R�3�yQ�GnZ �@�%����[SD]M_��*�Pt������s�Lv`Ƕ�jh�J��y9R�T��-=�;Ftȗ�j���i�e��%O
���h��m|[�ۮQ1D=�n���'�����ϟ���ș���b�$�2���8�U�=v�.B����_@�g�w��!�N๔�o-���[b	��ѱ�$!�9,$Dq����;ZbV��Ď�%�i��D���\%:�#��m��h]E�E����ψ�g�i;�&_�:�#��R��HRë��}��dF�8n�O����I5 0<���.�
�A�3n�o�B���:����mf��4LP���Μ٤��̷�����̄b��[�m~��GNF;GZ��Fs�ݱ����k��j�[9�^��ɝ�z$�4ŵ7ebw����J�C	�H���_��B��ok!���E�\�T�">C�EhL6/��* Z�x�R�O�0^�*�]l�Q�������~>>
�����G���X��P��sf�Es��dЈ�K�
�P�E���;'5���:��R�B��~�«��=�^��U����q,�qğ�7�Ī��N�1�S^߆hvs'󉭕[�����Tj
���M���yY>	��`�X�UϬ7�@z���P'|�r���t`�P�����;�z���^^��ȝ ��̰^o$�I�i>����^e����؛�E��J����ݚ���'\4ԕ0Dq.Ԣ�8p�.�t�?��c%>3�y���9l7!���Q�<K�Yz���"�����#�'Њ������wt�t���v�y��8t���'V(����ۃ���fP��ɏC1���D�����b�S����_��M��Ծ��c.�ڜ�_4E�2TJ��C���ݐT-7bz��Q-�hQR{;��bQ�P�:@@��OPE�2�a)��io�'���r�I@�ʔՎA(IO*�]D|[:]�^m�C�{r��F�� ���Mkg-�3����4�mw�!��J9ύg��Xy�v=P�	���(�hp�=Y��\��:R����׷�i#4��!��D��kPĳ|�d݀<Ԡ�>("V[�d��#��z��������������q�Qo�j>�;��iF����T	7�2�PjQ����m8���߇���sT�����=���%4��l3GTW�U0w)�w�;����e�SD�	<�/Pc�����F��Ij!��=�נhŞk���C�u��cK�t�R�wj]�t�H�EE�Q�N �
~;��ϣ�\�M]N���D��!��6\��ա�]��(�V�����(u�gs{]!!��s?d��{�� �K��Ӡ�҅?�؞iWA��@�R�;ޒ�7-���0٬�݇�Vv�M�7%��Ez���L���h��=�����h�
��h>Z#*��
�*?���_[f�ko���"4T�ӂ�[2�	��o.�!Ԏ��釆υW���U�_�r�7��Ih
���S���
�R���x_Qo��$4<��uP�j T!�1�B�
&[u�#�ҍ�&f�v�j�N�Q��kE�&v-H�y�L���<�>E�*�"��H{ītf�˾�'#�$-��g�w�sL��KՉ���U'z���fՕVHJ�e�u�X'9��O~�ñ�o�o�+���X��e����|+ȣ��u�cWe9`�	d-���rY\�j�cy��K�@N��_�S��Si�x�O��%��{�]d��&�����_4�UL�������JHc��	��}�Y���+a�/.s��N�:�%���O�ak���u?��۠���4�<8�2̰iGʺ�')$6�T�[�÷B��3��Z�ɉ��OK�P����Ax~K�f�#�����;ٓ��<E����}�[��	��*1dV'�I��t5��5�.'G͚�ܗ=�]�8Z@��(Qϻx�Y�J�d��jj�h���������IBq=(�����q4��������;�?^���g���cF���6�(��&!�Q2_4/f�����LT�f�8>�C�ey�p�<Jm��sC,K#l7�Ci��-���&':<��5��0u�!��������o�@�1}qP�f{_��2�-0q�#S�)zj����$B�fw�:�Wo-
Д��C6c��wt-
*oq��UVb �����X�8��x;vމ�F��ܴ���޴��,",y.�:s��?~�.\W���#�j�t͑��"�c9�@;4}<]Ú� y	c;�39Qȸ��V�5�8�U`��۶ob6�P��C8p��w� �f��x������o.���`3(	��}EA9 6?w���d ߕ9&�MՅڸ�s	�E���R��g^�B�)�*��d"� �r�}���f��\֟U$n3�({
3�t���`��B�v��6���M�U<����}��{��b2I��z�[+����/�����E���!���z�������U�/���o�A-�x��c�r���ˤ4K�v���Y6���5_(UP�W�_�`��b���E���/�E��p��ŵG-q�a��-���q�ϧ�N�<����6�
��a��d)�?��$��`? ꊎ�i�R@�ͭ������X�Ě-R�28� �?l=S���z
�u��H���{�8�"�
��<�U�w�'�2��@~�2@Kk������br+|w����AK�h�����l2ҺIROj�q�� �(_�2K�!�����J�v�21u<�&\��y$ZAz}GP��(/pܷ��\y*,K�g�-8js��wY�����j��D�D��U`�^����5�k(7��d�ZSe���T#g�LS����xn�2IlIr��Qó�kZ���.IIf�`�쥯��-~Ġ��V�LjW;៞��p�A�y����^��=�5�n��s�8��vh/~tC�{�{}轋��R�*�l���6��%�"Է�c�eED�ЖI�'��D:�yǑ�hs��c>�Ce� �?�r���)C��}Ls����0^`�8F�{C���D8��N����¾��F��K
�>�U�s�-��緬�P�S�����&a~D`�Hݑ~I}M��@
t��Ȉ��y��A�XS7�V�fQ~�j��(�Z�7U]Vq/L�k��vw8!_UJ$�Bv�{�-�Ţ�EiH��o�,):´�������#�>��;�C�+��q�#��KN��}�Qk
v���"�j&3�uߣ�,��R��?架⼡'ڧq����h�K���{�Q�'c������ǃD�$Lմ��w���G3l*%��N�Ҧ	d�Ȍ��d9c��u���7.�g��}�ʣ�_������e����z&��K�xFl�(�?w�Q4�CM&�Np����"2��o�|=��߮�����ۈ���~�1�P��3y�1U���/�e��>�Qz�g\LWy�ձ�N�Xhb���"�J��K�<HP��{q���'���Y��N���O��OJ�]1x�4���±�Ҿ:E� �����X5+.��d�H~�Μ/�F���b��<P��q��"�Fu����,4�ך�������>����:(��@��0�-#����e[�F�ۦ��\�O,��ٹ�3�)�kљ�~��.y��$�yzY�
���d�>*5amZ�*�����(i���49�@�\�����*F��{A����{��EҸ��-�g۟=^=�5x���f�$Oi@5Q��\Jόw��̶}U�"�g~��O�rFh0��)�2tL�_M��*fk��.�f���&�=t��SPKks�5�.O��2���.�i�i6�\�<wH�S"`/�퉟*e}/,�^�'ےi���9��Ȅ�I�4&�%�R�L�6��#2k����vq^�n���b�W .R���"	��O�V�����#q��V��0��i��/W�(^1Ɂ�K��"w��'�|��Т$1��V5d	M�������g�b�=��@ȼ�����jw׌�]`N�Ohs�xW�=ɧ���E[�'�8)���f�je�����j�{N�h��L���N)���P?�N���8��s0
T	O��
F���	�� �>��7��|�̽ M�"3��6ķ�/�dP�Hѳ.��R� BU�VȊ���)��Ǻ�b�{e���o5�n`c�	ؚ*S ;t��0�z�ѱZ_BE���"����r�=8T�L�t�蟁� "M+JΙ�<�	����_k3ܥ�p�H{	����vO����{1��Yz�&�fN�[�uo��x��џ7l�����y�0�\
4+g��(��8�#{���k��6k������n5���'����é��1��Z�4��%��S�sm�L���R=��1��d�ߘ���j�1��̾�>j�� jwA��[m�9�5�{Aف�x�/GT��m"*��U����r�JC@b���<V>Ae3�0��]3k)+Ӄ��g�W�?���ĝ���}�Q�+yAv���@Er?O��ʮ�v'f��*B 
�7��@C�ƴ��?����d1?���"���g(�lA�`j"����a�#�;�ߑ����c�j-�p�n�x��m�����]-���)��S���o鈗kA#�` ^>t\�`��V��rN~�`�"5rdP�D� ۠h�X�n>�0��겾{P��G=�4��4Щ��{Su�������Mґ :2es�t��.	$L��B�7`RE)���{y�l��;w�ۿ�'�.��Svy3J�G��� �������5HE�ǌ/����_h�z���+����B�5�U�[�?Z�T�x���Jp�7�HG@w������� >)����̶�ۉ�=gٍVa���z&�S�:��,JI�D�h�U�7�S���TT�����Kة���+���W�H��L����Y<����:�l� ���W`�/<oWRo�?,�����<���<h<�/��ӔD(\d<m��U:�u��x@{�>��y �SIj���A���;0��>��u�g�J ��>��$�u�97��x�!�w|*�o`�e���w������q���m�y�и��뼬��Һ���m�豓r	����&���E�m"��^�҆�4�$�y�	���Y�A0~�K�
����{����^[���i+32�*l����Ǯ���
�A>�b$�����4�\w���>��d��Y���O��Z��4# �,Zy�D���4$����61I7�X�JYȺ����c��\8��~�aM0E{oM�I�P7G��ʂ����*wJ4�[�����S[3�I&��K f����;�I��(�~���Spb ��k��vɈ�ut.�G���4�\�y0jn�G/0���p}�ņǉ����y��٘\�2B�Qu"�Yx��� �rR��ZE�D�oa����#Ŝ�q�k�F��՛��\1nj��*H<SPwC� ��_�S3�K`��hz�@���23[C�f���.8[��w�!&
�����?w1��r��:7�����27�BքUEf˒.��Q��#k{��0�c ��ŷ����ϖ/zL.�����>��^�O�Z_NIӧ�R �eos���� �&γ��H~��n���D'B/r���v90���x�Ze�~/�0݊�|v�/�]O��x>--<��N�JJ�l�����S3�&����ؿ��ɑ��.e�d$JH���r�Q���{u�L-+�&%�ky	��T�+|��Pu��MY ���u,�2SU�Ř��gt7�
k�н4��壘{@���S�y�p΂�_2�K*���̇�kF='��p����[�4:5Q!�=ҦVA �j�\�#��M}�>�Ab�Tʬ�p�X�偽�L!Om-����I��IKyS�5�n�%�L��5�>d��AQ�f��NS�b߲�g�D��x!���k�W��Pa�m���b���c��H�aF�_޳��ρ�x�pҌ7ҏ [?�> nP�v2�;� �M������ɲy\ͽ�"���U���jB6B5q���Cճ��-�������c�!8��յ�k������)І$Ӑ��4A!o4:�Ӛ��b(�Y��O�FE���
�p	��ga��w����L7K�l�u�b�;9"��o�ǿ�gS{]{X1F��B�+�����s|Fu���T3MQ|^թ��p�26�벍G����(�� ���:���
���Kʧ��� 7CzzhA9�j���/���rE���\M�M������w�2�l����.X��Ypݷ�}=�׷��t\EQ=bU�Q�MLS?���ǹv��&���L̶�§s٠��Y*!n��!�k�3�%��6���'	�`o���`���&�1�'�s�m/�y`X5�\���G1r�с9��ene�W��f��ޫ8�A�T���������cu�ɮ��N������G]r�~��j�rr�[�K.�8M̼��h��x��
�tl-�����<�;e����� ה+3T�5��9�cE��J�ɪ1�v���&���A�!1_3E��
٫p$�n��+j40�;���R+�_���R�G����l�:�=[웵�Yo�`y�KA��3\��a/vM��o��n����qIa�1���>�/'�R��8k��,%P2���By�:\��Jx��Ǯ�{"�a{η�����p�u�*lĮ����>�>�A�t�u�=y]�$*	#[��G�bzI]�^�Q�]*pL:�
�-�w��U�#�lC�'K��k�gս���`I���p�8Խ������,�c-��X�}Z�������zh^��-��!����"����aV0 �I�}��W&���9�\qS��F0��iDZ�zf�`�t	��	.a4��Q�NP�[�_3�m�j�Te�Z��7`�/8�ץ�^���H���"�"�K�XԞ�7�-�o�k��~|�ۘ�8�^�؎XY�4�7��40_/hhZYD��˖� �T�C�%<�Pj���9~�e�o����]�V-�%G�r�8� V����T�K�T<�X�5!�3ێ�0�%�x���$q#!H���iR?�Q|{��z� X�h��U����yk�� �o��6�F��*�>��S�(���������P$��"�I{ٝ��t6"d�֒������V8���P~����Z_������P�
|Deox��`Z]�����E�P���wʉ�v��}C �T�ˈ�?�<��l�N]�Z�N6(��(�ģ9�p����-��R]�\��g����t��S2D�ᄨŕ�li��q���l��Tb��^���j��N�C��>�e_�,� F���*��g2D���5R>W��z Q�PQ��j��U����N[�񡱜���L�:4_bƛ���&�?e���m�uQM���I�;�Ԭy��>�"��N���VQF��xk��+�C�3D�V>m�p�rB���D>QM���w~��f��u_��R�clS�g"5W�=9={�	�C+R���u|�i9}��Sq���@cW�d�y���pФ^a���5��	�z�ˢ�?*n84�bsw�iC<��.��탋1�%���&�VjqA�*j�uA��R��_ъΫL� ={�	b]�2��&�?�E�MgG�#�H4�!c�^H�Oh-��#~^aّt���-5X��V)����y^��7��5�&B���k�~ɄwXL4 ��+O7�D�tP�N�Y��������r�J@
���o3��b���v���u��N��=ȧ�4P���A�jڈ���S
����zq4�&��A<Wź�M�W@�;H �]5e�#���Ո�?���
�)�L*��'1��O[�Q�� ��kă8�ySν��?�yNE������vxc��R�y��������!���	,�W�y&1���h�	?�m�D������\��}�{���i�]n�2�`��+� ��
8��e�Au ��{$ɂ�6��/b�5X�Ur|��jL�⺱�ڻ��＿{�v� ��{45	1���1�,�G��ʙ��x�3�y�����W��"��/Jʀ�t�}rd��~��'o��_WY�$^��-%������Yqe�v��hǩ���.Hk&�XRfD��Ɉ����3�L0)��%�w8�`�(���n긭h���~�(���M�f�" �E�7K�:�|��	���Aj��q�
܎�
���o=o�{SP��i�0ܪ��O~�_q���S�`5�3
���6�GT	�ǔܘ���/�M	*���7j7+�/d�YxlvAa�.�\��;y����T��Q�:�敦�X[��f_�յ��<�~��^�M�qoU*��s:V�y��8i��X~��fEA=��\�q��j�R���3�	�Y���C�V�)��{a�wh�"�#BΓo�Pu����Ƞ��;��}�P�r�Jp�#��o�q�z��h��q��B�ߡ