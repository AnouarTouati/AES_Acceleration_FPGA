��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&Ű��=�b��vT6�4��L�b,	/,A��"⽰k��b�t�u�zU ���� /��QU�:�4��u�"�wP^��P෤����?|�q��[�A����6G'��Ð_��=|���Pm��&
V��u�6g9�"ۓ�WF����ԥ
��� ���6�0E�
u�����o�BA������9~���lU��WY�,�ڡ7�  tj����L�=�7���B�?MF�	�%���ކ5P���gi���O��!Ҁ�ؾ��U��ۿpb � �Cc�{K#�1��4n��`[�M�jTm����P��u��� ԻS�{�/�Q�xhW�
�%�Ñ�sv���ʷ�q�3�ێsqSi ��NS����:�n��LL�_�Y�_l1.�u��m���[�Z+��ޫ��(KoMO��Z�͟�h�N�
�.}����2�׺�MUg�ٿg�О���k�c%����S���ݟs�e~��vhB@*:>���nͻ;V�X��h;�_;�
�1���L���w7;������5�c�b'����a�Ŏ#�=B+w�cv�t�(Ӵ�L��,��gTW����>H$�o]6���?#��[�Z-���j�7pW�O)<a�g�֩���J�4�#Q���U9�I:շ�J�m�����̨k�!}��,��u���]�X{r#4>R]�ݘ�	��J�sq����,d�Jۅ(�Y�B��ẽ���k��NX���?�=�;tk�����6Z�'�$��o
?1c��J96&����Ƕ�A1�-�;�
-��9�U�5�&c���%�q9������	�u����|1�+�y��n�:O�nх�a�?�_+�#d/�%�Q�<6
_�m|(��gh^u�S=�T�����ޮ�zّ����/d�LCT6rNfҗ�	ۉ�[x�Rt�9B�6]Ȍ�@�_]Q⁎�	Y@��I!�1�,8{cڔ��G;^���j}([��c���0!k(�����%�e�}�;{'	�دG�V�8���V��/e�vQ�}P�~�+��aL�>.��	)�'��A�i��6d�ͅ�	����	;g�1���.u�����E����Tyf��,y��Ocڐ�����\��.(8�o+!5�)��S?�L�N!ĢZN����5H��K
L�c�ӓ})�	�V��a��tƁ����a=#�mK N�P)�@�x֩�� X�i>�"���yDj����|�\h&�X�.2Lx����m.ɝ��]����ݺv�Ii��fv�,�����<���FQ@�2�rY����F�gq��]��l;�/I��Kv5a--�b'��5']&h�6�0Q!������opd�-��;�z��C�)n�t�xG�=�E!�0ȅ����I��i�"��2�#	��"z)�̄�Y|;�c����"�{T�Q�)i�����O5s����&�t�b5/�ܓ s~Z�R���ت5�"G��8aE���4���W�(�8�9�g��7�S������/��|��P\#'_��`�^j�������;#����lww��t#
��BM���C�^`����7��(.*���������Q�rR��R�#2��� `�����Ҧp@�KNCh�`�|}bع\"�1����>zj��oMq�Z�4�A5%j��>HLSG��<�k�E�h��:y����<-�hU=��Al�y�r�)��m�v�4:�o��.P��+)&�1����l�Ol�|��p�R��p
�a3�ο]�Y��l�nV��`0F��I}�� 8���^M��1�.ۍ�]�lڜQ���lK���Z��ߢ#iH��'�� aZm�QEs��G@�%�#_�=׳U�8�Ĵ�?���u��S:�2X� #3̇�h�����%���O���ۦcRG� ����+�^*@6pr!`���|H_�Fޙ�^��1mv������-s.������E唘�{��Ty{�Sj��py]��Tsb+����b���>�IV�Ǫ�@p����� � ]G��`�����r��C�Rϭ���W�kdt�$��,$����>1f�G9ۉ`�_�xOS�!0 ��7ѽXKN�8�H�>�`J&���IK���j��үM��֚�}ɴF�f3������U�a��#P�J���h��crK��!���
��l�Hkd�.Ms4������ $�C�_�E@��uŀ�	�=̧ß��w�
�>KM��R��UX��|��Q�픹�\E��J�4�^q?�9�3����cLqey����љnm%�_(`m��%�׍5Q��J��/ajX30�l�;�b���)��	P�f�
Uz��D�G2	��*�P��7�k@J�6P�Z+M�r�k�j�g�RfI�=t�+�C��TF�鋂�^ȳ�R�T8�8���z<&��$7�rXf�\����Bo|9��!�Y�4�����y����.΂W'��@��Z~HM5y1�X�p���G���"��&TD5�߈K��[GWL����
��)�ܘai,��Jx�fkQܬ��)"�:�!�H [�s2��87�(�������fB����a��l'T�����(�r�;`#��~2is�x7�#R�\�N�ԜVou�N�,uK�d�з���ܤL�Q��:��X��w��?*-+�.$�;�r��Kŋ� ����[hOIU��<�$� Kl��j�p������\l\R��f��;�:�����d�G�A6.d��D�|���RT�I�M�9��dֵy~�I0v���kN+A%I�j����ٗ���Y�aS�!�ȸ�[�.�O	֝��>�E�Ѵ���@���Q�5ٝ����k�"�?�{C%L2��7�%�Zތ?�L�S��Hf�S��mM<��J�v�sR�GLPi�
n��))Wҩ��Ŝ��ͫ-ÇA���u����}h�*���s"�o�S���t����<K�t�4���Yp�X�?ZR�E�X�o���f"���cW{�q���Ǡ�S��lޮ�(����C����z-n;���0�ä�V"�t��
f�hD3y��aC%?P�4�?�0��'�1/S���w�Ҍ������E���P҈on�boDԞ,�%-`��r	��|�����\��sĜo��#9����E�U,�xƜ�L��2O��pN���8Y� �k~��)��s����d�#c浥�_�?�=9��� �w%79�W ������\a7�G�(���c�s�P�D ���N	�h��d[�|ۙъ�d����L+6b*ټ7�?(��p��%�XZD�	��0h�A�)���'
�p���4A����:�<ޖ^�m.2���~�O���������kai��xH���
Wc"9l�4|pX���ln]⌿��ƫ�`CG�k�QZ�H�~�f�n֠�q\�e�����`]eU���$�:����L���5뚓��F��{��Δ:z2�oV�=��~��g�_U)u��>o��q������W�B@�b�=E�;��!^7�U\E�WS�V(�,ԻR�t�f�I;�|ڿ�?�g)O���r��.�w�D��ҒƗ�\��p�M�H�+�\o�i:��cK=ݍ�J�H/~�����5d����$���g�Ԗ��`W�+�?��-�B({R����&Li*hr|��fq;4!��]�7T.�&{�f����u}-��-4��Y�r �LBF,�ߓ��l�X��@�{|#�c`�R�VtĮI�mk��Ř�B�g# os����ީ"�:��-��U~5��#�������7m�|>�r(V��i�SI�^B�UˊW�ٚ��4����4
r�ѭ�֙Qߒ�l���i�@D�>�j�cH[i��s�"�*���)�+[�$}�ՙ�z��X�Ó��\�j��YB4�Lٷ�XKf�X3 *V�RE��Mh!� �j���}J�������εlǝ⭉�"����+��g>�w�_��W��!]�����u�ұwc%}-E�a���E���J���:��/�L\z4e㱫���SX���{$o~l=v�k��Z��!����&�R]Yc����&�!��%+��D�΄��b�M�RЅٚ́���J���{�7�D��U�ȁgi�%��W��?�l`�B�b�5�<C��_J-
Y�y��nK��
�WT��_��\ ������'K��H0��e�]��5$<opw�8�|@���t4����b�j�N�����eI�v�4rp�E�xo�IpH�*GJ �A襊�L��G��Vm��Y��r
�!��K�t�E��"�\�����!'�Љ�x�I+�h����]�E>0��&����8��!��>�P9;޴� /l0��?����	=�� L+���Ԉ�G-y3z�M�y]���'|)*���V��GjVz�U�E9�=c���h��.v��e#"Jfd���`4��z�����ۻE�/�ۨ}k@W�r��\ך�ʨPtH'ɕ��B�
�H�`U|uF�c
�P}T�nG����V���(���2����k��:Jr�������JF�ݖq�`e�q��0+E[B�k0��kp
>O}9�z��f�5�i�)��b�+���3��,���80m�9B;bt-b���Tm�h@G�:8.C�F6��9%P0s���~�5h{�N�Êq���tuqdej� �ː�p7j�+��J��~�k�ػ~��9�|�3�ĲGO���<D-3w̒�#^��d n��z��DQ�.(�I��a�%���Q^;,��&s��H�p��i7��$�kɍZ�S�Gr�bq��hk(m�)�W����&�(k3�j���������7/[�A�&�b�U����mގ���0��tc���"U�-�xh�FE�p����ɪ�P���U>T�ڍ�EQ�nF~�|� <9Pӷ�^j�g�������G�n�� �h*�f,�#A W�&L(v5��m��E�3��{7���茊��3`P��
x�,׸r�L%s�� ��BƇ�	��g���-�f��euގ����iSJ[����YGD8������d|�l�Vh�̵�f.���:��E8f��eK�[ �y�4EȂ1e=���t_����zŪA֕�^Iz׌ӑ0�V�=���K��=8���O]ꑶ0��W��3D'�^`/��zРbw¸�b:8:릕���Q�̮;��B|n"��[���H?��U�Q��a�&ß9��A�`�Ն>[���Tʅ�W ��5�&y2>U�O	p/`߱mN��	 ��r�ż�S�\�%�3��c`6O����A�_�5�I�7�a���������3 ߂Bx�=���J>�Q�ؾ���GP��G��i��P�ёr�Z1�'��&y��Y���b���oo�H��@\C3��w�}��o��l]��ʅ|?c���W�Q�xK4�x��(��ʔ��A�����Y�@=���C�%pm4���7��Y�����/C7�̦�VD���38�U��r���W�q��ɕ&,a�������<e5�r�0�f=��b�z$�1�Wu��ʪ�1�ׂd���Y� �bU�����;�h��f/��h|��NϿ����ςɽ�*�6�qn�E�G`2ow�O�^N��i7� ~�/����ck���>�;���4�?�
�D#�|y/��K�٩�q�K+gV�L	}ZcY�?y;,ń4��J�!�Xx�����0r���;837�����3]��\��q��`�:s%?�����{,a��,PK}����8קdkI��:���}����#MXs��X����#���������C��O��m�.@���`?��mA.�Œg#���bB�q^�q���ބ�H5�Fҽ�SKuOJ����lo�v!*��
c�s-WD��=Q ŚL��
u��ۥ6y����Y�<9]����J��I������	g�
i!��5K��_��%�'	�T�X��G��&��QH����6���\�6��L�{��h*�{���)�d�>�n�N�UM��� Δb���� +V6��>���M�ɔ&w��GWn�ia_��_������?��]��&�$`E����NQ���Rnu��b3B9:t�X�Vɍ���٠�y�����g}v�h����e/f$�AOu��P߾!׃����r{�L��e=m�n2ҟٞmZ�,�>��
�QV�6���;?��aa�ҕ`>�B��S
Z��9X��t5]�@�U|���]#xct0��2j/>��7+/���(e��^�⭖}6MB�E���5���^n���}j���0xKwQ6��i�^{�WfGn��v)���������
��d�S�>|�"�)C�B�S�l�P�@�V�)`�0�m4|��Y���L��τs<[��<���2����c;HK3�γ;H$wH����z~V�p�짫m�?
�^�G��t���Eˑ�}K\e�����6n$ ֛f9E�~$�����d������q� ���P܍j(`g�<�95ʒ#9��q���¶�MN�x�s��O�Z���_/�n�X!Q	Z^2�.�7y���5�/�Tx2�k���A/��-m�Sˠm��H<$��]�@&���s�ѤBԺxEV`rLQ2�Sp�խ���2#"��^�!�]�+�VyQi��xt����q�>o2&��=�"�hBF��=���嗝ڎ�'~`��P}-�sV�ŅQ�͘�š/'b8�{�P�i��`���h��lJr���66=	
H�ݾ�ao�ˡs�);_ýV �_��֒D8x�+��t��6�Q?镰�n�CS�%�h��{̩�UW��,���L��.�ͨ���f3qt?����Ŵ��>6B�	R|Q��c�(s70�5�;P[~��
��fg�~�'"_��y|�E�a9�Vd,����t��a���]$)"�����Tzj��X\|�G�V��Id�g�Jp4������ƠRF����&h�t-(��Ɏ>� �y�+���T��~陦����j�(ڥ%~:/�J��M
z밼;���n�#ٸ'5w	4B�V�5{8�)x�ͱ΢M���p���tU�.��������yNvY{��J�=�K���ШO$�u�"�v�b�`X��l^���
����|�P�/��1|�-��u`�_"~����S���lw L��y\�3����'��e��ʋ�1������g�o;6�q���}��J���Aw��j��+�XXG=�e`��kX�+�H����/�}�pH�;:���M#(������c���`(�N�W�'��ci�k�~�\�[�O��A0����!x^�/A�S����]��ln�q��QD=�狨|�ꨐ�� H�l�o��Pg��ђ饍0���mF%��Qk�Al��S&
�(U�{����&�Ū�V>�ZH�r�V.�;Jj�%�ǘ�1����oW(� �8�!��o��Ȗ��ma�U�r;��t�-˸O����gm�m�@��d�F!�݃��]j)��f��g��eg�]���}:���_ t�f#�W��;[���������q�+��(^��{�/C�Uh�I�-��Pm�cÿȮ
m�@��$-�#ݞo��{���}+�8>���\��w�fR��NS�ճ��ϙ.[2�7�'����]�k��8T�WEUkYU�iJ���ApU&ߑRT-�7*�a�|�P���!6/滽� {�!���{���.h�<��%�%u���g�������Rm��:��\���@a�����l���3&�X�mV�}��FΪu�>���}=݃�p�߽`�m�Q�~G�}r��u�hnc�RKg�^�Dü;�Z.H�[��>+yK�gчV������}�-�W���SV���GP�Զ�1�
� ������N�5�:��X�%O�a;�$kA�p3��m%^���Z�d��C����&�כ�39h�U��W�>PP�� B��l�������G��;�3�/�����N��V{)�R����erk�f� ��W�t�2} �j���4�ݔ�0���h�K����z���?��4���m���Y��^m�t�.�ɶ���R�^b��Fث���`��"'?�%ugbv+���p�A��q���[��a5�ҚhW���/���� ,J��۶t��C%qE��_WDp�,�"V���=ͅ�Hz�.J6��8�\�|1N�zI���u�O=���,Ke=S[�f�`�L��y&/Q1���C�0��xUz{@���r(��>>G�v�-k�+n~,q�O�u�+ޭ@Y�j�P\�t)�e�R'#�dT�e���|�#&��@���~���)}�H�e:RNM��6ɿ�ؚ�
#=@�f��d����ɺ��|a�1S�z/�C
���c@�E΁�W�I�7��',m��N����9V��+����#J

��-���}���l��q���Q�Zy�o����=�D��-�M�#�?�U�CS>1��R|�Cx�H���#�Z�0ԯ�����"��y��X"�YO�������?`��3��Z������^ᾈ(	��@y6����aˢ�U���q��Ǯ��} Ƣ<	N���@�[H�+�� �Eu̜G!�tPVwHݺL����K����L������S�*'*���c&&RzYQ΃I#=`?�A�Z($e'�;��Dͭ�7��e0ǧM#�9?%#�,��sa�0?&m^�QHB+�(��d*)�2Xq�No���f�
�	X��.2|�d)ɇΩ�e4mf�D2®M��G���$o	��
T*)Y�
�
%���:�q�0!���+���D>bKXH��BM�6�W-�H��p�Q��$������Iq�$ߦ�"���p0�d������Bu��6���#�H��t�s+� �qO�G��X�DG7���6�g��"3&��qH��z��қ��tؖ���X�-�Ӹ���0����K8��F^	��gHb���HpM�	���L�ǿ��ڢ��ܹ��璿��O�]Z�ڄ������]��5��c��7�nAU	�0�����AE��̟w�vxYcXg��n��h���w����Ѳ�ŬF��eT�>V}�+�9�0�Hr���C�e0����E�P������r	a�º�,ϝ_H�6$�=YD�Io��ܔ�	�\h���)kD^�|w0�R�N�ы���z��C%��/������	�0=�3��O���N�2����Y�i��#]=���ȁ5�<8�����d=]�g%��hY��[�]^� fW�W/L��d�j�-��i����MH���a�hC�E���$�&�Ud{��4ؠ~R�����@����1u�#'�|&zY�oCɭ��]̵����|�͖��#ALy���Z�y�7�`A�Cn���/=�ov/B=}�=�w�� ��0�)�2�I�gʞ��u��K����)�"y�/w�ph�1�Ut8;M�u�}�,���ȃ��!�ݜ�N��L	Q9�E�B����i=�M��L�����_�ܵ���Eg_^]|3U�{����-A���d�z	w�%�ZE��?A�"}�{�Q�ȫ�嶵�\,s������������Z�E���gkj$Y���(�!�V���`�ڊ�l��s�S}����~Ƅ#O8�b
�Ҫ�U����q��If�j��3�2��7��{v���Dj����jҒ���P-6U�Eo�A���/F.�$���(u� �f�o�	d=H�:�i?X䛓��Y���f���*`�b�p�q�
�\<k?�?�6���M@��9)��,k�r�mO��c��" h��r�*$�皌�J/D3���@�b%m#���
!d�����[��$��[#�K~n�Qߥ�7`Qw��e]K$0�uAK��"�����e��)E�1J]���/�&��!p'��3x��;V8(��(m��ۯw,N�ww��#8b�y�ʝ�#17�>�, �b�$����I6p�
?z���
����:8F�$G�1��uL�2$�kJ7����^���	G�T�+���V�p��#P��P}J�L��gX���v-9]b�!�o�QH�.�X�$�?��كb�Z,��^��>��W��Y�
PT����2D�Tf_��pmT��{᫖K��O�����;����V� �"���b���گ�<�K��I�M5H�Dg�����i�q-�����e�lJbaӺ��e��U��ŐL���O��!���zO�w�M��c�t�:_���+C֕CD���v���HF��B��	��YХ	�=^����QIʬi޲x}��&���B� H�)�D�I���1D\��K��q
=�ˣ��^�T�2���wNB��}���W�Y|W����(����7[@X+��eXVܵK�m��J�}��@����T-��Kʢ�hQ\/(nay�?�j��b���1t �87����-R����ln8K�*XR+��ͽg��7�	���?r�y0���K�*�[�ۤ�x����m2���T�2Ԕ� ��ɠ��0}S޶�%e�aޚ���k�S%�mX}�=�����m�E�.=���3��ɿ�|"�3j6y�e'���l.L/x��O���Z���f�)�xs!,Qпy��a!=��1�UgC�'�J�FR0u7�K�,V4�S`ؐ�f`������D�&x6�v	��'A=\�aY�xV�p4|����5�P�`Zգ3�촏��ݼ�-S.:�܍Gqf@IpRL;<�dJ#�}���a�J��{�R���<�.Y@��!D �iee�v�-_Z����!�U�% ����r
������Y���:�BX�c�y�#DR聋2¼�ϧ�W;�x`I+ �5��Ä��s�h!ԇr�EQ�x�ߏ�p���;�������»<#(]y9����2�3S���Ha�Тt3ZƏ>x�~8'ʋj�TL�~q��L��jw�&�jdq4�<5ఒc+Y(;0��/|��}���t����>:M�ͱ���gڒ�l�<`Nr=�k��Q9�b�3P%d�v�"C�Z�U�cZ����Y}]ӦC����e"����lи�\*�W�p�5��>4j3 8��<��C~Eސ���̼��C,R	�߆�q�Iq�iW^�+2�(�0��<�³�_ )ڻ7��[N>���\��ؚ��U�uY�G���s�V��������� ��F��}&2����f���`꾠Cw��"��K�ۼ���)-��:�%���X�M_.�R"�"L�_�m�B;c�Mٗ�Ҍ|� ÐLU,i���JaB,,�T@�m��	��kMC�ګ|b���qjs������f��OF13Ϸ��e�Q�|�qx�3�*�e`j^T�$?��Ua�m��6���{8��՗���t�i���d�D�T����	��W��q��$Y��H�V��2O�ξ�. ��O�npB��*( XLn�S:����#���ǭ8�ۧh����jj�0�q�%2 9��().��k�wY~�����C���:�nJY��G���a~g�VL�
J�`���^�VC"�����3V�N�- ̻�6��_{ ����K3�=��Vc�W��+.HK�]sgnۮ��vj ���D��lnm�>.�:��R��}E�#y�tq�'�7(�QZ��蔗��P�W��w�N���>�!��c�qF��C���P�U�=�c�r�E�H��	��U�dG'�F�)������4H ��Q�[�:����6������k�^�,����m�p�me��֒���V�o�P8gQ'F8UL/+�=kI����m�/�3.Pq�R�ۢ;�n�W�@l��Y��TBM?�s�J����9	k����8Y?���7��#��� ���!�F���k�X�ޗ�Y�R��w��{x����*+�p�KK��v�H���dq{�eWX�� 4�`�B��ԭ��4��h#⢽�a�K��Ƽ�g�L��%�S�>�Ej�j���f�O�r�1���#�zSٯ�E��!��О�p?�ɳ��s4��f%��l�+�샮��^ݗ�1�p��U��F����~z� �տ�/:�}�0+��3O$۞�3U��M,���C��F�ɜ�!ꨅ�FN��� V���,0^f�v�F�^
�b��(Xc��7mj'�.CL��٬��h"(Į����=rZ����:�2�7`�y�N�r'ħ�g���]E�h� �U*�rh�k���^Avu��`e0��r\!��h�N�Y7[r�u߼ބy��7����8���.���p�@\D��]�S�v�(���3,P�I�J)A#	�YA��[dW�8����Ń��8,-x=�:�@��>&Q2�2�L=D>=�:��Hw�p�����^�#M�0��=ʬ��D�r��A�'�-ʵ�mƮ��#~%<�|�a0#��7d�*�&�O�.�S<���{Kw<]
���\�I��^�3��_�Od����Wo�v�$A�y�wI�+�?LrFy�z˳����2�'�����#%�r�)v���JN55�`#9�����pz7�A/����\�a��N�,�Ԯ����*���:X[��F��3�!L�w´!�^�mơ��i��j�V�yN�ǰ�{���H�+��7��$����8���|��s��x� "{�����7�մX�Bї�'�kay3Ĩ�2,��3i�l� ��_�wY7�i���d��^g=A�0L���E`F������F����|�-n&��bIM��h�y�|d��r��$�CW�qoq�S��#����JZ�	E6������u�é�̝q__�NE��4��Jx�F�G�������g��
Ӵ�Ǧ%YE���ھ�A�vr�n�ָS��񅙗�ן�������;��0�s!wK}��w[9�(�ֆb��i^Ȧ��e�S8�'z�5o3ŝKlt�5-�/�	')E���E��w�yal3�ȶm����K6����"�Ф�Z��l��ѫ��3d\8�;}�X�f�C���qe���0*����:l��;a>d�b����_z��`�+��Vb֮�hK�V ��.bbo{�-gR$����Q8���w�.��C
e�p�Y|���'����$u��ADVkN)�����u�ZMrh�'{"���R���b�tv�JrDe�¿���1�8yZ]���O�H��	M�G4Hl���sμ/����8��xT��,1��hw^u�h�/f�A�=��$4w�\c���(U�5�-����;'�ض��F�:���'�؟p����jC����]h�F5�k�T���5D�h��A%�~n�R�a�+�b���6��`�!�hF�q{�R}FM��^�1��\Fw��!�vw:k� K3�����)�y�w<�B)��m��G*=�C 6�݁^�� �j�J�rTo�����w��� �o#9��+kI�e�U���y���.J�N��M�`��YQ�R��a��b=��7����z1�Q~q�ח+w�d_�Ń���Qa��r�Z�V�x�7�"0�E���Y���&��=0��3�r��a͢��/~#�
�f�'�|�8i�V���0cY����Y\�u|��шє�{�曺���Z���oM���D%F�qJP�*��,�s<6�|\t?�x��;t�Z6�Ra��K�>#�"7B���҇�o$ٓ�}i̧��l�b�ɥ)1��n�h<
�2��"������M!��-u-����[X���^���6;�qf�ԣ���Q�8�*%���.ЦyQ��� �@����>[8,10���A�
0�L�g./���`�y�s��M��z���c��58�M�K�ȴ��Z&�>��;o������M�
[�VhI�PU��[f=Z�r�����Z\�R�����Dx9eO.d%�͕v�����E��V峤$�h`�-F�;)#�r+�?��t�9���>2���b��ڍ �i��pDY�sƺ�����l����(�3^Čc^���p���'T��sq+���i��2�����N�\ue�\�UZ\[�WJ^-���k}'��@r��W�z��L�`/��.c ��;J��D9z���P�g�j]*��f.v�!����6��z�?��=g�{K�	W[������Ho�R!��-�Ღ�h��M��)9FVV�^��7������x��e�ܤ����zGD�d&8��S��%�j�L�/�����F�)��<�@���C!X�70�������:e���v�[|R(t�I`KS#]��&��ɢݔN��=2ێ}���8n�L��F�̵ر�	S;���-:���,�W�������E���u��C����SE+H��~�g\ � *�����l����PD�:K|������ڴ?�j�u�E0uL4,sC��3�Ѵ�9�����f��|ѹ�Ȋ����E
��r�z�4u�_dT�{��7��A8�L���W��C0x�a���V�}G� tm���7Aeܣ�O���2��7�DY®X^�.�;HO��QI��Zh�����|;:	�Jf�������I!lw3˵>����p)^�[�˵+S�����i��'�r�,G���+�pĭ�qk�wx�6�=��*�����`VJ+!�g»*FX�"-��Œ������
`�s�%��nO߄��8tm��H�����ݑ�Z���t�������c�h�{��Y���#QK�~.�o��vKz�~$�de����<S>��4�8��-��d�ҡk�6	3x&1�^��Wq(��@Jc<) �n�l��>@����ϟ��`���?ʌ��/��#l��86�_�{��	xKPX��z���R�|��'~������WE�f
�	s�P��`d�Gr����|��	5��q#�u?�J���
����*R�%���l�jz��1ώH��0_*c%�퍡%Lo���
��T=,�uVU�"�G�v�����W;��W @�mIQ��ϝM��̲�mZ���`�������N�zй����=ŗt�čڀ�H����"�a��,�{�{`W4�R=�tp%��2"�2X�oy���)/űf��w~d,�����,��.��ط�I��2�=�!O/�[�;�B8��:����=
5<R�-y�	�q�S.8q���]�+�1�v(�^X�Q*U�'<����_��65[����,��)6?8�� �������c����>2E;�0-�� 89�<vB�G����,�����t���K�X�C�E��ۣ�j���{kҴ�
mY�c�؇���O�Џѽ���R�ߍ0�شBV\[��O^�M���Ia��y�֠�4��.�3����� �o�d��	�3h�5�}��s0^��=�*�θ��E��B������N��riP�<	�X˅W453ͪƿyё�wU���%���?r�����ؤV��][�=�|B ���j�)�|!FX#v�Z¨	Rʎa��"Z)^���3��$ʦ���V#!E�#ő㨽EcE��g�^Sߎ��D2;r�QP��>�%I-���5�$[����2^��gPTx�Ǧi��5¾[�;	S` p%��T��-���.�f�پ���#�`�q1��=�ˆ��/��֬��VO�VO�gy���.���y+�F��V�o�ITxg���'LȺ
����I����*��M�A�$��p�2Y8brbca��k�N�{Z�iN�b:�s��*�kj���o)������������G?�����q�����؆��΁W�j�������䱟�����<7��PWYo�)�+�R�|���_7U�8ہ*�8a�*�I���i��ܠ���dm*����#���x~�
	�߃\��r�끉���N7��z�����p<`����v�Ym�h;�TY�o
Ã�M~D�@f-��
�ߐ�7Eù�O�*��۔��OH
��t��zIa��N���;e[*$�nudo0&���&�����n�0^�Sr����i�H��u"�5I�O�?���������0��>����f�[����NC��S�ޠ���=��h�{o�������P/�ιz׃ęuA2��Kyo��PT�H��㛄�U	4[t8c�6��t�+�LT!ٖ^Q�8_prq���t�0p��.�9���uƸR��(��9Vp�TC x�gB[���1��=�,�ġ9����zw =0�=x�;�4(A�9�H��I26t?;�	��Y
�QMc49��!���m����T��mp3�ȓ�-���Ta���i��DxXH��M��	�k��W�d�1��w^������"�1����D�-o�B��<m�њ�����)�NX��4A�y��O�7/��-�t�2��n���`�vF��g?�6e��#4L�d�Nd2N�ׯ�rh�RPi�x3uPf��x�[�Ӌ"����g�þ��Y�bR�^ �q|닻����7�[��qY�=r�N�����Ţf�f�(S�@'J�] �n�幁��!��Pqf�;�P��0<�����Y��M��)�c���X@��;�q��r?c��O�/ʨ	������'�s~�,�~��t�����1��9g�@���v��>��
�6O@����}YN����|�'�{wl@T��r%~�U��V�,�8�!$ݯ�H��8��a8�����vI�Ԑ���?�}���SrzPg̋��@���ۨ) �F�A�v�^8����܏e矎�=i�����a�"\��6wB�{I�
�3K�]6��c�e��x��kj���GV�k����!�E�o���[Dh����wёMg�n��Pf9���UI�\��q� �_O��k3{?�FC@Bn%%͵fA����e1�Ӓ����,"�m�m%�Y1�Z/@`־/��oTd�wd�d4���U�w�'N��a�a[�o8d�ܴ��j�U��9�g�M��^�Կ�tq�g=A��7� 9H�����Q��
���C_;�E6�Ӕ�{5����k�WvT��uw PX��ScRb3������:S�{<�7�"��m����]RLxmD�)yO�* ��4іɞ�E�.��uʟ�P>0@���a\] �U���C��G���3q2�Ҵ���~��Y�����	��f6k���H.nh��̒ۅ���`"�r�����'+ƫ��K7�E7a-�r�#������1c��FB��~���qC�F���2��I�bJa�pj�ٺ�RF�j��YK��J�l&�p|�i`�#X���ĸM��b[v�~囤 �9�Y�B��j,j]�5���鹸�n��݄=�9h|HB��(���V�)2T=4��3��wZ�C�AK�&Z���q��?=�S�ˋ�[Zz��ܺTȩ���7�An��Y4m�Y��&�	V���I�`_k�>!��q��6�;]DG9|+[�j8㟴"��D���#�}��Te)pa���f&x��}! )/C� �I��؀D�/�+�3l�����V ��7�X9%x�ʗC�!�W~���� � �8���z e�ø����pvѾ}`ՕVnD�R#���Tvoݸxs¹.�n1}"�FKf�}��+@�3�*�M�O�r`��M��
#���a�H��h�����,2��J��F"��`#�.Cu��f�D��[Xa�?���{i1;�θet���5���8���J��J�w�o��a��D�g�Yg��_\B�D)�]�P���2��Q�\������� ��=��o#b��nO����z�xK �gY�Ys���vt_�T1�u�7���/��I���f�
�~]#v��q�#��3�-��u�(x�W/��:�en�Q�������Ӥ@O����ݐc���Y:׷�c�S����Q�l����τޖ:ͣ���D��ʫ����$l�"z��M�]r�ʤQ|*lt:����鞠�Z�6����]�H�g(�Y/���+q�/�I�3���0��U�o��G��~��a�';�����u@s��a�{_��N�z4k�Y����V���kF����}C�Щ�j� �E�n?��z��F#Hi?�sw��	Uu�	Ѩ�n&�sAF7�h���ߵ�l��2�R ��g��F�`����ğ+�dZ�u4W�ˏ�J���ۧ-GC�=��3g*��y�7렝3S�O|��[�]KcV�Ϯ�2�����w v?�qWJY�������hJ��Je���-1����A�D[�� E��0�ƪf�E����*��9�3��Kk�v	6�U����q��(���V
ˊ���	�*�+�0.O���ӳQ��[�_�d�Y'a����w'�HsSJ��8���ʞ	tx��8��z�묡��e�89��,��:By�����l������4����2�aK�il^,���ե]c�°��ֱ�rWR�yR�Af9��M�l�U��Fp��?����E�=ٌ�C��f�����	鼭�&�Sqk���z"7-#�� �݅E��4q� �����9W�r��F�Ҽ�?�"2�%9��ۻ��1B�>f��<4�<ߤ�w4�˔'�9�4�/S.g�$ݏ��0A
C	o �īW�e�eNӣ���8��]�R���杴}�b���U	&�'x�3����V.lP��c�a
�=2��茎�خ̀�Թ=[��]�+������f�c��#8#�&�РB��x
�x��?,���.�U�˂ΰ	��5��[Jt�1��g^AF�s�w�ĥ��̹�~mr�Eެ�0ҡ>� ��u���]�f���-?q�k0��U
�z�Jc�E��(�S�b�!�j(uqJ+��xc�^��BВ6Q��I��X�|g��o ��F�/����߲:�	>��Im��N�Cg��F)J�͘��e/�YIÁJ�d*⏊PQR4�ӳ�e]p����@$W'���*,!2��S�,��ilm���d�y���hh؆~�1[��V��|��0�|�ĄK�N���B��d��nh2.;׉^�VW������U�%_,�q;�#e,L����+"\���6v���\0���|��"us�88�D�ȟ(�+#�֟�ӯ@I��i܆:\����6A��Tl,��b��ފW������f�R�Pyv黨�jS��^-�i2U�h3�dܓB~�3Wm0&A�]�����J=�2w#���j��^��-���`�Q��v�Z��Ʊ|~���5�H)��#TZab�NsM�78��%��R��'��� �؟�T�.K�F{�EF|��H�/�}��	�K�b�Jh��B,���@�R�M鷞������> �kP�-�
�繄Y�I�ׯǔ�Vr�^���<%�},x�"�JRм"����t5�{���ϩC"�f��b�7W�W��8L�u�L�u��r��X��)Y^K�2��Q�:��׊�e�;��:*"�l�pK�'���K�=�OAe��Nf֢ ��7ہ��>M�rc&�P��!ź�y���Tm;%�� K�	��}���E�h%�gp�W�|W%��Z�H��s3�3'�W3ɡ k��~µ��J��g��LUÒ8��B�N�\ ���ϼ�j�����/?9b��q��L��9Ƀ$Ϫ���k�:e���+����
����E&u�?�U����