��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&B/��O*ISO94�8��ٷvXC�!^�%=�UarX@l���[=U/��-3�/0��6�%�e�dF�(.���W���d��1׼6�^1�V_�1j�D�eC�KE���+%��~2A�P^���8\��7����d^ ;}�{~Ȣ��4Hm�.x N��Rs��L�`t���(�o��D7V��o�X�PŠ�7j���(
S;pb�r��[�k"��R���
`ٖ��dW5��E,߆p��yc]��)�
�κ�p�^��FP	��R/tw,VCO�� ���7~����A�����u����GȪ�P8j'���r��E��$x�G�-�~�A��6ֺ?����0im��k��X�~z«c7#�����6w3_ļ�P�u���cK3�����Z^�x|��ɛ�S��iD$���Z�:&vEI��}��$�>�ij�m/Ǝ�
�Est����IV����7�\�]`�f�B����l�ʌB��pOCT~껄���*YD��N��Eq{���I�)�{c�8�D���5������b�Ҟ&�!�a,�J��j�0���E~�G�`��Z� 9��3ΝY�g`=���n�KK�� T�=Y�T����t�N4s�l�jB�(��W^��պ�܄%��5Oʴ�a��(��x��u.9����SDsdpi �K�dםH���Q�Fũ!;�$WcT={�N�:����X�ܶ�^���K=���"���8��U�3������i8h �mm����.��&���|�SCQ%�]Y9�.�(�����8���h�;�s7�z�$��	�wႤ�Ce�>0��/oZ���������{E��5�E��T�a��4��a:�B�Ϻw�ulu&�]|K�≠�i�
w��)�a�ۇ�17�6����\�߶s�_(�b@��ty�V�y_˻�	��2Ы-S���SX�¨�G��"�H0EVX�f�I(�2,�#��n3P�eD}7���YشI���w!������V��U�a�UP��J�m�	��Pօ;󆦡�z�GFK�5'��JQ|#N�ʭ[��os��+	jC/H��=��qU}j l$��=�x$㌽\�9��G_��D�:�����T�<:��+��F�B�\�ʙJ��q��i�����7u�x@�`��q=%��p�t�@1��:�ԑ�"�X]��FlS�D�X2�ۚ�m&3�;�z�]ǫ��5����t�XʄuE'��7���3?�C�X�G/r0RWDre��xWo�TP��*h9ՈQ�6FU��p ��g׃�����4�w���[��?g�X"����{aMW�麕����D���S�m�� 3�X��]c����j��ت
yS�eMSޭ�U��p=�"�ﭺ����䃅&���?Ζia!p���,�)ue�RED?�������3®�K�XB�Y���w�Q�^��:�#�%��7��FS������'�����؟&��X[4ֹ��P��~����<Q�<!���=AW��y��;���c��6�s�GڨU�9l4���o&�к�����#���{���J�3�X��2�i�2w'Fg�o�\$D,h�t!`�w�W���z�o�Q��*���^�L}X��'Ԙ���3���f
� n���`�.��kKw��J���:�h�?�	��9��p˻;:"�bSo"ڎ��k	>��+7�4I�"��P<ڌEc2��ڪ��bˊ��;��e(5�O����/&rd��pz��7�t��ѽ�?��Q�Iqőq`�����.Ɇ�|�S-Fe`_P��}�����r`�H�$�ڏ�����M��X����v�?�����i�"�⢆��Ӟ^Jj�9K,�ߜ N�IU�����L�)<�
n����N����`Q�$��qf�g�Z�GE��<�V�Qv��?�W������=Ǧ:ig�N��Y#�rn:�#��4LNh��T���	��G�� ����_�`�vY��`�a�&��� ��������;����I/���*UtoT�_�A@�_��E]RN��У��%n���CN�6E.�u9�P_�p��R�ŧO���h-�jԜG��4A�v�L�(�`#I$��z�����/%��q�VI���vB�bJ���ͽ	\;��)��W6�-���ҘXI��.*�xY�~��}\��Q�8[�u�V����Y�yX�,}/oko����Z.�-q,4����>"��`������(&h�3���Yν�]��j[��T4Y�����/�F�1�b��dV�䴐 *}�E;��z��0nu� �'�Ix+������X�'�F_����F�tc�k�Mt�o�,k��u.d��УooaoAI�����+F4EV_���M������ ��*ؠ�5癆�� ��Ѧ.�!�irڕ�����SH��7hԎ�P�s:WJ��0b�L:Wyg�󾟔���c�Uh�cM� ��Ջ�-���=�� ��z��$��4�]�a��r�>G9,�"$����jܖ�tz�?aY '"��VްaC��U�_YA�S�����k6OFô����������J��{O��1��[~bl%�	U�o/�3�y����E�蕚?44G		.o�0/�W�(۔�)�pߋ|"Q�xL��J�C�`����R�x������C��O�$�s��QM�Q�E�Z��ik;�ɰ8�'��Bp�]q|���/�Z����s.��ų�=�R��E�X�L��O5
��Nx�))'�
e�#�F_���G�iݧr`8xB{8H1@zL�����҂���^�F���D�멍��6���)M�8�z7[/��:�3F�u�3x�|M���Gz'$�E,)��ކ�3�A9|v�{�GT� ��ŕ!Ahx-���g�ޑy� �m�#h��,��C�*"SkȈ ��[�O�I���߱6S������H��O�wWy���9V{�#��Y��#�����;����ƚ�(~���Ve�y�ť���D�]�I�aD0�;h����X|g�DE���sk���~)?6� %����+�ΦQ�GåS�+��>�rۘ4�Yv���oא�7>'�^�bZh\�9��#��UER�1+�k���
ūG�=�$�1"0�S��є4�WE��/5uL/;�
�g�Y}�}�qB�hb��r�={����MoC��k��~�t�6Љ���k 5�u��q(�ǖr����A��#������R` ��OLN��T9*�v�w��2�Z1Qi�0��6�S�H�"�0�
S���t�XԴ]��x�H۟����z�&k^D�!l�� �V��:��ZӶ'l�~lo2O}�0N?l]���ipD�פv�>���t;����d6-���4[
�i����UQ
�	�����sC	JZdܠ��=˽	��Mu���7�O�����������2�K ����]s����a�1m�"�J`��(F����Ce���-+���	��jӶ�N�(��@Y^��d�*wc#�	�)�p�����l��0�3��H��>��v+� :�P�+-.���S7�TN�V�c�)Ć�%��e��#���N�Aۑ�Ѿ"e���db���k�C�
�sy�X��U&���n�$�IT���؏Z���di9V�!�c΁�9CϠ	R�%ѓ��p ��n�oS���MJ�(��,p�9}L�Z�A�8?���p�G��:Aq�ߕR}إ(1�d�M�_ѝ��
 �bM�~���	��|��p� 1���2T��I�q'2W&b֚��g`Y�i�g@
�xa�;����) ���k����@[���>�pM�w���bA��f���v5�ح���N�� �e���d\��3���L�J���Y����nO����m�x��VŘ���u���޳����؅(țJ����k'��n@2�)�#h��[���U�ҙA,�P^�6t1c��G�fJ�c��v�X֋���/�1��so΋�S��'x���0"�CZs��s���k�;B.oO��){�T�a�G���(.b�U=vk�\�����,�̰`+l�.�`�`��`nL(�	K��)Z��1$��Q �k��҂����*���+���X[�dǅe��T�A���[�e��ڐ����:k�0��*�p�����K"?����/-;�/G�xX98��$������p�"�N��^9j�<1!���6?~ţ�l`4'm�5N�u;��拈��w��Ҡ��5Q��G;xw��!CsB������֘4�����AI���n#�#�O2�f
���\*���:��c�Y�P/ￊ�,���,.��2�����^kM[>�&��\5�fl�6���~�	+>_���FaL|ԏ�U����8u�A����@�8�Ҷ�!ρUv�-��t�(:�*��P�8�.! ��ڈ�`;�$�3(����3�P+���~QC�����(~�b�p�r�b/t�W$�$��_/Ot3�H��in��r�KxԊ= �$Z�T��8Ź�����v�m$�C��(v(G�D���4v��mښ}5i[�ӵ�
;�Z�}�kQw�j�bu�"��I�J]{��zO���^}m�@����%'I-'�r8��O��j�Xڋ#��ޥ\�i���Ck��W����"jF�Yac�4�*D��WL� ����Ǒ<0��ݰ��%�#�� N���j�	��)H���\wT��>���&��G�u>KΒ�1����0ȥ9S���;ݔ��_�w�|���{�+M�33�-�h�c�~���.Lgb:�9�u��6��3���������T�@*>��`ʢƉ �z�� lI:h#i�%�����Tأ�'��y/���b�6)��[��VrSi�JK���%�.~_O�m�D^m�/�B���A�Uɭ9�rJ����qi���`>�1=�˘��w)4h�*9�dk��8��A^Q����E�#q��Cn��Uu�V�O�3�f�"�Y�K�mX��߾�!2 ��%���3�z݌g/����}��)  ��	���Zb�˭Ϗ�t��0����&��Gˁ��x2��2
k�*/r�%�?G(~3C]T�HaD�g,"=%��q0I� ���Z����3���t�Y%�D�����{ff�˃��p�s{iŰ6^���7�j�P���F�c���&>3;��!E!FĊ��>��������d(�%��E �Z�Mѥ�K��'Z�+�c��[�״XXx���UOhu��o�'�.�� H��]���l�Y���~Y�ҍ��bc7ۗ�u��~^��3}�#!�G�}�������Ƨ_J��[:�Ò�M���*r�9|U�=�${"�9�t�r��잺k�~�E=s�,&�������ٯ����b�:��^deKˋh��`��|Ӛ��)�V�5%J��� �H�q�.*��B0���iu\7��1� �'w���g'?���P7'�9#�^���O�efjϭ�7~՚>�8w+T`q����Ue��AE�Q	���o`�Q�j�����Y�0%��͸q�S(��(v8��Le!�Y�[&N�j���4ؑW8æ�xST���_Ĭ!�0���="9�t1��.|RB[l�b<9_��_䋱�Q*.ʥ��ّ����:LB�P$w��&c�|��>����q%d̤�7�\l���V��$�ǉˊp�_�!�o��ho.P{G����M,�UB������0��)��B�#1����v�ޕN�l�����s����x##0:J�h�6Ł�#Q�W�&����=�#,%�ޑ�h�E¹	X/���.�1���C#�}�<٘u{�E�D����FQ��;2-��j���'����|��t2?f�ĭ�"&ч��[��Q/WXqq�i�}�2���,�J�
�F��3�M�(� D�ߥ����cu����!�M�����>���bo��a��pEҪ4�fc�pA#�xJ+`��Xh�P�A��I7ۂ�ﰨ�P�w�i����	87 I�)�0#V7�&E��:�s�=T Z�2*-��D�t)�e����]�X��x�Ќ�<�o]PP�&�4{�K���+���O��fs�n}��7\�$�$��A;&\���	i�G�L����j�9''l����Nw~�K5N ��Y5��ɦ������;C���_ �m��j>���pX�ŉ�®�h��: �(�O�˳�"�y��v�¢����d�Z�ܳ�?U?W�����Rv���ʆ���X{��|5�o3C��c>��k����)��fZ���߼1"i��,1_�u�`�5�\g���A�R��� U?~����r�\u�'��Z�u���M��\�f���i�s��U��(FɁ5�Z�oΔ��n��1��Q�;���(&p�����m�t��yytc+�B�{!��Pi�Bs���\�r+�ȴ\Ѻ�yHxh��(�f͸º�v�Ϥ��������p�y�d�ï}>gU|����؟�#J��� c{/�*y����K�@�6P~j;�FKO�^I����v�6��Ԃ8�Kw���\���2��O���W��qo�Z�Wg����|sk��F���K��8�\���ak+πǝ�F7���Q��l;�X�"܀Z�t���|����ph2��5��	4Lۡ����ؤ�X�{�_R��H���`g�*�z�72&��u�]a�"B�ǽ�3;{3���q�?#��s/�;76����H�Ji��V��#w����Y\Tw^�6�zg���@nhX�2�YZ�g����G���> �ݻ���)I̮~��K�9�!٨�U����ِ�Ȼ�C\Z����Z���s5�!}/���%�;�,�cB[��}Vb��`�RR ��.��"��uc�w�[鱭S}����z.�P��J/���V�x#.�r�����S+��F�&�V;�Zҋ�*����Z�����U}0&��j����Z2> ���>�ٔ{Y%q7�&y�44Qq���%V+����m�3)uD��{�j�笤q)��2�@��(ޝ.a+��K�|�-\3�����p��]I;N�g��웼}'��_���\�>W��k���]兕��k�� ���E춁>��=t�o5���D�k�;,2�R��iqS��`Q��NH�4L߲J�ip��e�輵����z��A��9d�q�`ϭ��}�
�R}��P	����׻��N�4�S��K���K�G��A�H�a �oz6Mz��[8=�no�\��Ĳ���׎�x���x��͑��}�}o#_��qy{V:��y[|@���OϏ����<FI�;`�x��Mu�ߧyk��[I� Kf���ni��1aEdO�D�Z=S�������/ڊ@����s��${ϗ�q]5->�m�(�UT�,F���i(	%������d��n�f�L�̉#z�\����˼�	Xj�F�1��xB����?9�{���`g��9ԭ��K�����pI�y���ivd�N�9�c�8�D�%��ʪ�TQ�K���:H�p�^W /ʑ�����q?}$ċ�&���RQ,�u�����j�/W�)�����)u\`�h�`�۽;�#&���\�$f�	��&M�3�l�k��I=�I���ߖF���~���#b�U�A�om4��P>��ś"�����ձ�����~������DP�o��)��w�l��(^Ŧǰ6�$���Q����W���1�I��(t��<	l\m�,�c~c ]��[d�Gxl4�e_('I����,�r%�t���n���� 7"Bznޚ��Ɂ��ك����Q�s��ytw��-i3�]Н�N��X�:���Wʄą��Ki�E�C٭� �Q�J��Q�|�D�����wk�C���Y�v��!�ձI�CPu�`���3�]�.�7���ZY�G4����A���rϑ\]yauI�3�`0� �x��v�V}Щ!�IW���9�z��[6"��ƢfI�Mi�B����/�'1J��ޞ�E��On�LD�sT����gB����BA���Αդq�cz�+W�:LkD~�߮�ґa+`��B<��e�׍��)d)yWՓ�s�����XL� @5��8⏼�e����	�:�8�B΅/�|8M頊�F��G'������C���j������B"F&g'���>)���*qW;∽�R!E��<���t��+I�Y1J>m` &[-x�]�����
���kǀ���gT�lif���	����r�Ts�a�B	��-����Ա�7	>��}f8�����np�O@���=��1��"/��/�1�����I7����R�����=�����ǂ�2�\`H``J�:��0aq��D����1\S[�Y��T�/��X�{y��}o5S�^�Hh;R�D���j�����(�h��H����O�"���Y���8����Kuݼ��+ ���h�>�4=v��&��eB������c�ҋ@,���n�k�4��,B�����4("�k̗�2?`"�ʵ�P ]Y��C˕>��	���ş�kn8IA�s%�u�����[1�Ĵ�Wѭ[ڇ��EP%X���Y���fG?q�_��{��jU{R� &��ةŔ�$��ѸA���Wp*{mG�Aכ�̽��gS��w]�k?�R�8V�fuRv��Z|��G6l��P0���C[V����hC���v2Vd�&zbM�<��u�㜬�N9�e*�"�=[��s�IȀ ѿ� ߏ
O=������qbp�(���9#�W��"Ų#hD�ID�`�(���$�σj�y!P~�k�̭Ճ��}���2�>R��_l�}��>�̛��_?��d7<H�t��͉ ��ݪ���	'/��wC�a��;�gw-&ߛCӣ��0������.\J�[����[�����oJ��d�:j�߃�n�
AO�F DyhG f�"�m���w�+�{����]�()O�;�34Q��e��~;>�i��@'�@`�X/�8@xt��ܨ��������!b:�_����1��{��7L$/2�"����z	��ܸW���E��d��B��tG2Z�5�9���]��XX_�a�
���ey1U^9��z:��tUe<������G;�/�W��z�H���,�J�/�@�cm����[`�3�V��Y�?s���xfVh��\�� ����>T���9`m-�G
�Lb���hi�(	�P�{���0߷�~W ��n��fd�����r�9�#S�ǩ�L�)�W�"�+���T)*d	=�����DuӔ.5-� ���sg�Ji���Y�U~����N��B�&��A��:��y]ơfVl�?���]O�֗-��c|�w	�4s;׀+n!�J�8pG�vC��S��t6&�w������ ���'Q�7. ���JO;%k/aƟ/`/�����Y���,䐃#�V�`w[q����g��`�ɤ�����uO}ѝ�b�}�c���Xgk��QĮ��xӬ��|sZ���c!}�f�A)P=�����ܠ������j�m�����Y��;5ѐ�a%��Y��9$�GB�b��o#���;�z�p�и���,H�u���Έ�$���Д߼��y�ޠ��*�a=�Q3D��r�Z�xԘ~,u��{b� ���!>IC����ۧi�:r\��_�*��XW˩�_+�YNZ�|K9��x�d�u��W��j���O�,�H����d��|xM�K-w�K�ɜj/� ��*@�e��94f(�T��bE3T
Jf���d�ӫ)�T���ǃ3�FC�˭q>�"ְ
&sV��y��Nz��V�E��+�_�	����^����K�g��H����Ƣw�=��%G7R�o�m������H��2�+]� \,��N���r���?|�5m��D1�%�0�|�	m	75,N����Yft&���K�@j��z�VBu_�%�/�p��vw�U���,�Gb��\<��k�p#;j�N�c:ӕ���K ��aA���N9K'�Bh���@g�#aP����*�r���,uU`ٳДg�jO��4K�Y/���G8��q�mV�O"�Y�py�S��7�����qɀd����F~��ĎHa�����+�h��	��$��"TY1�H��}c w~E5�bP�g+j&�&y�Z�XQx�g<�a,�D�r?=������C�t(��c��+R*pz�X���S���M�Ʋ��^�����:^��La���?`��{]����%{��\ �r{��@O�_uғ7 �S���������Qc]M��d�D�����ၻ�o��6��!F���v���U����eGi�a�?�D�ǶN��dr�&�\���kG�R{��O�hev�1�7�,khy����FK�U���5��-uW&�/�5����ԅ��{)p��Gw8>L�v����DɵwU�HT���RjR�oN�ɦ�P�x��)��*��{�ĥ��X*`k�l���G�C�7gz�Q^�Q���
�V�T�e���&-�7o�@zN)[$ܙMůC��^�U�ؤ����ߋ���혡w��o*��YKFfQ|������Uu�>����'�'�#^ ��	Gf�`�y^�Ĺ�f����j�Z�ﾐ?R���t�h��7��[�#ֿ(Td�
�5�մ'�b�li;d��U�~D������;%�`�6�P�����!��:�!0�'��XZ+6���[�wxP�+#�t�J�*�A{��#�3���^;��|��j�z�B�C��nE�3���9�<C���LU���&���>���IBL�\��W����%V1����M��+�%���.ՙQq?��s�چ�-�l���6�����S,�C(J�M��WXIx,Q�bP$�&�V<���ۡ�����4���Ek����ؓ�hFɢ+m@�l&ʞmDY��?v�_�5�'��6���;��+����<bbft��9�5��}#��ں���ۘU��'*1w�
X��qS�����KYd}J�M�(��Z�˵�&���^� �P�.��H;/�Q����	pOx���o�����BU3�������������@��?����&� Q�݄�)�po��I��n0����^Q뙥�Py
Zj�z�8Sq�YچD�;���S�y�����?���x����~7����E����4�ar�!�@�mĺ�
պݡ�bIx2���9��JH)��葨��G�E����S�V��wBhg���]x����i�-ܭ�K/�%)��b�5�`Ӎ��{��V�ޡ�����v̳­E'��zE�I��h>�H-�n�)�P[=s�tj���\���q�T��O��U�a� �q_xO�s���Cy?�u	Z�ek�W���$X4�'�E7M�������f�$]9T���!�.���n\{0�
�\m������a/ :�w⏹�t�s�0�,t��ޫY:)\�^�O�ԓA5�팆O+��|󇼄n���n��t������&�8��u��u0���(�h2[0S�R�:�k�$N��|����d9�����{ը��`�Jh�YnD
�=k���� ��&۝b�+�c�<W�%��T&��'xO!��xq�E��3��7 �)ߤ���`�_��d�j[�7��Bu�z��V�������h�w&���Z���ml�͎�b�C�!��|�����>�ʺ�ޔ*y�����β���ݾpP�R���RJ8�����T���.tCX7�B8K��{����癅9'�m��CY�Vyb��ً��%��y>��P�d�>�m*BA�#�� ��u���]���YH�2�m�@'$���!~���i����]�ವ�H�ߋv��ϥ����϶���%>s�ih��w��ީ�=�L�3f �`�jI��1�$7آ���s�#:���G�-�.K�.'!m;������麒�q�#����D��%�<�) �1�sqE�A�嗁��nkf�i��A�#��FLAE���tі�zYn���n���}��^%S�����uA����UU�rI�ܹ�'j��Z�{|}1��V�	$Q5Q�L̈́0@}C�0 �3�]� oKOR�8uU�QEvJ���{�l7X���2��(_j�lo�.$��,�N���$0�로��WƱ%D^��)t�#�wRA�����nb��ٕ2��@T�=)�l_X��Ǧ=o�x,����T��C�/��4���"�O}��3�{��do����7�����0�uT�N#bw^�j%X�}'��	��{�wJ�d;�k��#<+�u�����K���&	: