��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P����^�*��H��ʖ��Ũ��@��9n}�蕬��25�}��J\s�S1�+���@�2	����X�fC[^�QXv�0zID�?ͬn��=�W�7`���n�،��k���.`�	J�ބ6W����Uo���?xVC'K
RI�=.Ą!&��g�>��w���I����؛�횞����֢D�u��� �X���w�Q���b ��'߀�K�����Ό�V ��B��<Q�ڠ?�� E2�vw~䫕EG���_,{b�>��k�	��(SĂ�3^r�S���K�`��8��BA�ɖ(
�&��iWJ��v���^a�/��:��3x>�@��,�̻��#9��e�KV�>,®p�M�e���$�y$!�(�.��90�����Ƶֹ�M)�S��6�ϡ�h�N#��+��`�N�	���
I�D�^�ަa���1�/u��'��ʀX�,��H��ރq�>�$������|'�st��	�z��t�hrgj��j�\Pj��"����3w��MA�5c�\�	Iq�����@%����;SͮĜ��*��� �����-��]���{#ERHWE5O�c'
dB�=�)����; V��	�`C�$k顑����-�	�je�c�X�u�+�y��mc��>�;l��kk(=�AK����4���_�
U�d��UTw�/\L�%ŉM��vR��_-�1'cyjY�kI�,P4��'���,J�U���:'v���9H�N�FQ���b�!��w,֪��!0}�(�3�eс*{~}O�!IV�|���	b]�	��}���ٌؚ���9+��c�*J�_��U,��}�6����z�d���|���n���~L�_Ӻ��:�j$�S�=�$�*g�I����gn����E����O�'����+-��*�to]��Q�6�/:[�����Ҿ(fo����$q7�@�'�k��N-��Dśj�B4�д!���'�R�����Ԫ6+���;�(���y];0�Alʡ��ť��(�Re�a��BωK���������Mȧ� ��{��h5)�,g��̌��s݆�&`d��̊X!d���a"������Mw�ܾ����ك�X�N!�#1��¥���3x���V�I3�?���d�v���$��?�� ��%��+z�����4��:{@�p� ��aE�:�&!" 7?AMب�I���_,Е=�
�/�?����#������/g��]��$��������,.l�Jz�.�;�������:�|�82)3��饨\L�r��v|V.Y-�K�O��TU'h�M< o�6�t9C���?~R&�/i�"�j��rd���;UܭA��QNW��«��,k�L9�\R�@0����=H?M��w�F
K6{{q��OT�U��3�F��)~�*h�8�I�0k�x䦍2HMD��,�ܾ���MD��;�f8A�J������R��(���z�<ـ&@��b�܊3�Ͽz4&dZ�aۣ��NBBZh�>_�}�nf�x9�h?䏞��%��Kx�:N�zH��'�(���c��Ԉc��-���� $��⟬���6N�T��l�,u�@S����^�R�Q}�#���M=���{�&e �2��b%���JK_�ϓ�P� ^����D��!�\����2?������}�����|Isq�hg3�M�X|
��KxW�QC!GW���ņH3s5�K�Mڄ����H'�\A��O�"�U\��00Ǵ6����cά� �L�5 .��lg�:H��w��`��7і��4d�a=�yP�!kX��3�X����8�>sX'�����һ��4�j��1�ye6*uda>�-M	��T-��#|�R/�_��%�Რڹ����C�-��zPp��a�P��]n�q���˞A\H.�	��[��b� 
� [��	�"M���Z��\P,�;X@��#��t��79�TN�&E���Oi���s۠itCA�:52f��S�j=9`E��/y2���� �k}n;B�G^0<��B&�^�.�v��W����8W���O�St����_���'�s��z�\�g��9
��,�*�9V�ܑ8m���Q*V���ʶ8tQ�8?i��H�]dqn�����Zdm��J*O�(W�Oq7Ŝ�s�#ް���"b�裡�M�~����a�M���(aV���Ȗ{�����W��6^���\S��:�@}ZtШl2
~�i��NN����:�͗�o�n�͐������.J"��f��+�h�/���-��]TD$�4�$�w������X<�S��a�@e%��FӍD`�I��Y��w�Xcx �s���?Yҙ����<Mr�QʘS�3�"��mW��]b�f��8N�l����C�и��U��`F�x�Y���l!�(����%��wAv������e&��R�*����q���	$����2H��n�`�Ivs{��� �A��D�y1>�sc����y�	�[(z"�A���<�~<��}��,r�ؖɭ�@<�a��4~T~�sl0�%�� Z�����+o�
vű#�@�*���[#%�p#���#F�V�ԣ��o���(�a�:����,盠����Pu`��q�q60�Zi)'H��Fe0{c.._���]6lZ��)Fs�l[^'�",t��AC�cU��ɇ���Wi�֑Z\Y�B��E��J�(��і�p�\x@�I��	`�(ʺ�R���/v`/ؒT	B{���b�A�B�R���*��fLb��K�نE��M�[Gj�u��}���Ah�m@�G'DS���5�ȭ�]��7U��!�m�?���XA��ʠ˫���������vsv��Cn����)i���>K&3��*g E�` Ԉ��8V��{�_:ck�L�ܘ�ژ'L�ڝq8fߊ��Mq���f�M9���
B<�0=���,,d�bu�TU���O�A95(�4#���UJ�ϵ�q����3�µt�wB�1]�߾ݿA:��	_���u&��7B2³A����Tr���8����Z�TJa� �@�� ,�������M�끌P�(�۪��kԛS5gW. a����N��
�¯����z���ج�r���&��/�'袀f �f�<�q���,�?��Ќ/�����Q�BAFP:�4��S�%)���	�(�;�N�V�{40[q��:�;N^j��D�����n�X{S?�ٗ��H^��/�v���q�2s����ͫ�;���iT��U0OLwt���4�3P�o0�@���{�b=�ڐ	�b�n����6Į�(�*�ÁX5[%}BC�%���F�o�"�`��/�"�M��M������>�XZ�6�n��+y��N�K��?�QW[�:�fv�zM����_a�7�'0�?��V�u
5m�mg{�g���.���`��}"�܎�4��=O�;􇘿V5L��[�h0����(��S{�3��l�l��8�!�����`�e�
�؟�d����aD�I	R�$�3��d��rwǂ��U|�D�-G�Ӈ��}�=��b�P}�Z��W�s���13t<2�����bn>��F��	�Pu{��P"�~.+��Tc!�?#���/�c�|R��Hc����ymV�^�?�R�Ф��!�:�������Ӏ��~.�َ��Z��tv��@!���|n�lѥG�W��u�+�	]��@P�@!MiKS+j�����t�o�G��6�V+��p��FI�.NsoF&���8^q�a�P�»x���U�����yf���HB� 9+E�(d����&��>��mq�	�}T���ռ�j�g�j͆OXw�;��	�������w����Ɗ�C��Vϐ���wK�M����YL�r�'f�(��U��{Gb�P���e�� ���q�{�P�0��i/_�.gOOe
����Fz�\���<CK�L/�s��iޖm?9�è�vhXq���0>=1��p��{�&"��1'�12&9ʬ��f�yK9���`��B��?I��R?��0V��K�C���[�)xD��ͮ�DC��n�da��ڜ��|� �_�q�Կ~�r�
&$`�Ts�_�V0G�k��/����at���T6r���@�"���3� \���	���QP�����OVS�/��6 3��{-�>����u�N��ů3n^��ZyM�e��U�c�{v�܅�s+��U.)�x�F��Ķ2Z>u�
���l=��F&υ� R=���c��W�g���1K4k5O��)jq^���*N���G�n�En���׿��My�=��7Ap6�:,�������_H�R¿[��7�dQXQ��+���"{~�̻Ww�z����M�L��+C�Rp�ZV�"C:{���}B�����0!���t ᲺC������H��«^���B)|�8T!���.�sh���F� ӇEeڏ��d��tm/*���oC���S�g������K���,�DI�^d<��X���7J���C�� t%x��Q�7y7(�ބN�Ñ���rQ|�V����	`��[��S�a�'�v���άͶ�A%����&S�3���cM���!w|)�EL/�bd0"���Lm���ݛ�d�|w���p0��m��P��gb`��&����L����;I���a���O�}ˮ��$�l�t!�]+�0\F��rݙ�cq��`E���z8��:gYD�
Y�B���'�[�<�[��l�S�ɒ����d����N������K�m{�]����\̡�ue��+_?��uJ�pȬ���yZ�� r=e�VՆ�^D4�I��V��R� �n�[M�-���������@]�(ch�UdK�ɓ"�&����c �G#5ɥ�{��� տ�B�uEc}<g�;nL&��O�n}��/z�8x��;-Q�#�g|���.���<�y�RN�!<4����)`�j7<����x�y�b;�����Y���U��2g�q��)�z�Sy?�\������y�2�9�K�/�?+Xj^��Q�r��\�Ww��9K�ྫ���^#N�}P&��y� !�DP/�xG�؜Rؖ����?ұ�^@+]rpvXeP�}�( Y��l0qu?�(�PN�=dѪ�7�z��x̔�7<m*�Ow���UT�gm���o"oϒ����Ւ�5v����#s�/�y�jmz-.�#$'�3r��Ml �����Yq��Ue��ꕺΈ�����[��k���R�e�����{0��V�P���}�xE4�q?�t�G����K
�<���J ��D]�.L�WH�z�T����9��S��5���݆���d;���G��v$�x�3A��,R��Kχӈ:�?k�[g:	B���ʒ9����J�5!fr[�9w� h�g���b@Tz{�J�}ЍwfK,�64k���gݘ�Sp��s9�����}�E)Ǚ����B�����X�,�>CiĦ�w�5�]{ڷM>�6�l�<A�Z2qc�cc<����K5^;�O����Dݖ/��L���B7�MOUS��Q�!��l�]�U)R����33�&�N$͘���"}nv|]#�{3$x�[j]���v`�7���J� ��C�J�K'�Do����|�`���~����Ǘ{b&r��	C}��PWU�U�ү�.FDJD+��б����lz@��f)�sm�|�ܼ�cC-�!Q�iG�>�'����ٌ��8��m�������8�g��4D+#�W螵T��&�#{�B���C��"1����1p�����8RLW���Lȟ���w~�o�<�S]H��m�)��{�y�o���h����D-�T���=�o�z@����I��W�H��]�`��S�%j�7�^mq�[�)T)����%of�"ؔ��2��I����[�=Kv�'=R�goE[����K���	)?i��� �i�cN3������.Z����n��)�e��w�����p�2��!f1lQ�=t�V�����x"�[���� `�O���]Ԅ6Wp֋
IP!tB���] &��T�dY�����lgO��c<��1�.�]�X��bȤ�w�b�yn�>��k�h ���mhY~PVk������
-�~;����jT(jω�����._]"@��ƭ!�݆)`��15x��x��F���"u��x�Z���=���q)]1����+����!�~ʁ���:+�����sِ.
! 3�.�����iktHN9�k�$qhOr]���t�NC������3.��l��/F�ڈ��mwL��њ\��@.����s����|�i�q������E�f�<"O��H/��Z��ϋ�E��2O�G�mྎ����-@Mj]Mao�ŤI�q���yo�D&�;nf��W�����c�|��v��EMP�T	��{��3��M����{&����WAFZ�"1��{�^$��l�Fa�,�<cTF8 �ޡ����5yAUgo#�ɯ^�!J�K� Oi��y�5�M���DQ>��#u_��jw�q����_glPϞ�ŗ�5��(rU�X�wyZ��b�	k^��x�$Xo�߄,���[u[|���#���P���6�x�N����[ i&�ਾ��ZS�m���z�2���u�;�<��&!���$��D+VY��D/&�K�h�0�x.0�^�5y��@�4"[�Z��W�y�r޶ �O�"P�C:[��8ZDض�&�S�s��|&��[@Ffeߥ�9e�Oג����_�PlT��ɼ���A������b�d�tk�/�<���������eY���t5Jh��5ۄ��x7Z'���)���=��W6�Qh|�^�$`��s����넝ҐPj�4�G�}iH.i`�>�4�*4�6?I�W�S�1�?����A�h��5�P�N�N����JV"uY�-�s��i�y�2:+F$�HI��U:��q�'wa�7�v����z�*&�S�m���49cUW6K��S�P�����>_���G+�ko+5d�`a&��VNhC�o�bR�S�z�|!툌�:����w��Y�+��w�٘V��;d�瘋
��i�ظf~����K����jש��[�z^:\`n�h��%�n��ߴ���7��x�6�V$��,��H����L�J�B�	�0.E�7���]�E�O�%<�S;މu� ��p�?]H���0x6�?�Y��݂�-�.��E%�ʩ8,��G���z�|�tY)ߒ��{�S'�D�D{�~�@�/�qB�[�y�ݝ>ͭ{�qn�d5$��t\2�t!,юm�����J�^y�5�O�0����-Wʀ$Ɨ�l>�H��&"*���$1:�����������D����%�A]�`Xg��<nB��,M�C-$����d���0�x��o�x���Ĵ�ZZ�hN3j%����V/|�@����
__��9E��
����"򍹴��ш�+'q�������P�}�~]x>�|�I�f#Cwhs~7 ��w������9u!R���@;���!��"F�� �O�����|�9͑��mm�e
ןa )����ޑ����ĝ���!;��*x,3��GBZ��D�4�������e�KcU%
*K�KuW�B��4�F�������Qvƺx�k~�_�=`�~UDQ�t7gv��X���8S{����m���|R�i���M5�E���hK�NX4��:�[�$�m�v�g_�?8xĥ�O�,��;�;�Z�?廀J���!�zM/egr/���=*��覛@�Y���yz��G�iG���U:-����*�׫$��3���'���P����B�`F��I�m����C�L�i:W3�Ū\���D��o�~�F��((g��sE����g+yۍj�ȳ��]ZU����j������K������,<"h���\*bU����(��L�)�&*o�PF�V�^�8�l#%z�->�,K���K�D�(�;$� v���.���
r��JZ��_u�y�}0m6*�ac%nt��n�9t�Bϭ�@$ʝ�Ć�q�������	�@����щ�ѪlA��I��撪��]Ԥ��9I&X���<��t�;9���f�Yy�
�c�S�Q#�S�	��o��W~!�s�arU�w�\q�p�x`��������2� �Y�t���%Nn��ve�v�ǭ�}Z���ꃌz��Ժ��ƪ��$��~A0��.�h�M����@��!C@n�1�Ֆc�fZ����4�&�O�F���z��v6<�)t��tv��(�J=��T���b��Э�ۙI/��u�׸�a��zSNXh���4V���_�n:��\�öZ1�Ծ��c�F�{�Ї;�HA���J�x�.�-���WZW]��0���D���^'����[Y�N1� 	d�ۊrC�����=��c(��:�N�Ħ^�-7��֏>��"e�����Č1�����X��UHY��9\��{���Li��W�gX4r�?̯�i娘�|�������|������^.��ߢ���fsQe�o"��;<�xW���?�]�/T����w���+������4;�1�s�Ӧ��qp�/�zt��vv�w�j1����r��=
H���5�iŤ!��ܘ�"����&7�{w{
|���Fh.�ɥb�0(�T�+���ʙ-�(�m�qc�',����p��uS��e���H�%����L��j���DJU'��=�f��	��5B��{�
�ɹ��.�E�U�#61�"
�K���MȜ@�^�j�y�M4(���G���ݵ�Nx͂bW^O�=vp|���bhq�j�w�5E��΅�Z�SE�bK���|J�!T�&a���k&�n3��9(�\�6# ��,�)�/p��ǎs�Q(t�F,�Z:����'�y6�H8;K��Q������mD��<C��q��@Ĝ�[o�fP*�f��xw&껣�`�d���T�~������S��GGU�8�He��]Q=��=��l��K�Q�᷏l*���?1���S5�Ev��06����lz �C���b@��2ks�k�v�F���D�ǔmC�1/�FF���D{&���.��9/��fL�� (� ��Na���E5Y�
�5{��H�	La�Zc+g*W� �
8O�v�>�=�d��g�`\��+l�Dx���]� }*��W�²@��/��by.[u���i��&]n�>d[3�SK~]�t�����_��t��x�� ?�uO��o���0�x���vD_C0ץƑ���E��+ݛ�����X~��������I��[<gF��4�X�����wy4�<��l�  CP��Z<�j�p��!7�d|�&|�Ú׉���g[PKm'�A��hz�d��g'�TR��l&J����TX������uk-[�,�C��`���7PK/S�I=����_/�@ρ ĻK�"��mu��í %�;e�
g��>㥞���ǒ�G�ɉ���#N���W�".�e ��g:3ǅ��a�;@�v�<��s/����	2�/uLL HpӇ��vn�S��)���6�7ScXu��#2����ɺ ���LF���ub�P:l�?,��kM�E��.`̘�=�����U��l����<���k�\�U�$��MW�@�b��z�F��LCmv����w��q;�=(�xOS(��mN�ڨ9�S�R؃mn�O�x_�� ��(� +C�/�/F{�}ER���ଡ}�I��i�Yq����s0Cn-���kot���d�- #88X��\�*,~>�3S_��2H�[Ǆ�$������v�d�խ1"���~�*6�ᛤ�ћ��
H���8��J����;���ٌ9����O�ժ�f{9u+y���1~�����n`^_X���T�5�AzY^�dnK]���u��A�$��8�����s-�w �4[��d�"��	��V���(�;�qi8K�\��}�~o�X���I6uJ8�$��NxQ��V&ȟĀ�����i�����Yr�Lb����$9��w�
�͍������m�fL5�݁�����b�N�������n0���A����\����5��L��ٿ���<a$@����) +�X.� �9mq��3{�*/�2�H��K��:#�b�e!�2��&���l����$����!=D�{+~�֢�k����$b-�;�?�nܸ����z5��]�(�4��8�[�Y`Ճ^�)�R���=���-��4�ؠ�)b�u�B-���动�*5�^G=Z��!h\�;S��u��L-95�w��M��;�F��7�̲�|�ؗ.rP+�GOI�=�D��g��Vl�*H��Ti�M��Q�f+���1��k0�OX�i-2�'�J�� �ؖ�_���f�������]��(��0M�)Q���l= =MX˲iw�b&�F�K�:�:�&��uJL���U�(�(y3��5�����WM����=罄:�M�N���g(��3�R���M������ ��Df��!��%�ū6q_CT�t�\-�kk�J�Ʀ�@a�v7���a+�|�:�O�[�w���i`�!�������\v*�"��e"!��(�AK]�05��/�G��3�z2��
K�ڊx(��aw��ӫ��������D�̈́ �%3E���;r�>��K��Q��F䡞�sݰ�p�&�1��+JpIaB��@����Nd�"\@��6�A�f��9�)��m��!�#�!��3Er
:~xy_�4$J<G`o�㋓Y��FV������h/=������L�>���ca L�ggk�-Oon�T�יB��)����N�I5ʡg��b;<�%�%�A5_��QX̴H5:r����l/@a�*�$rv&6ػ0^ٕf,��V�秅E]�Dܴv�m���:M�`0���B��7�Q/�����09���.��u&_� �9u{��\��d�~ɮ��OPN�7v�
7���vҼv
}�<�[ў27�zT�s�����K��1�~��}��O�8"c�� ���5�Y�@�D�
�aF�1��P=�*t�TsϘn���W�rk��F$U�u�8H�Vu�L���O�Oml4}�I��2�唌��5�_{�X��m���U�{?��7v;��AJ�d.�neEy�\S�h���y>k4�
٤LC��K�WA{���4B��eߵ��Ϲ1�#y�S󘞯ߏ�h# �Ǚ���Vΰd�쵳8��o�uK~���r�O'����#S�k�]�%M)!cI�L�͗��W�D��i'��p���)�_���������o/V�JHvɶ]�~�B�4OA��6�(`�G�"B5���⸵��������m�7�މȐ�퐭�}-<�[_u{��� �}E�'���o�j���]]��ibf�yS{K�|ɴڪ}�+��gR�W,q�1�SpZ��D���<�Idt�{X�}T�2b��}����85�P�Q��6��J��
e?��@A��ח�ο�� ו^���r
�n���H�3�[5�iD��BE���)9ͫ�rk�=��b�k���0��K�@����K/*�O�YƮ�eCÉ��X�2�
��;~'q�;г�̕ʔ�;�N/�ȏ��:N��mH,<�7���<}��E�Z�d]�9MH9H�*dd��MOY������A�!*��$��T��O���t�F�����qM.z�X��]�Pkl�,ryC�"-|D�`*4�C��_&�	1�؄G^U�q���E�B�_�<U�x��Piq7N5$�&�,�]C4�Z6��W��
���C�
��T�1�䠪O#��8�.�9��\L*[�WD�P��Dˡ k*U�+֤
�.��)�E5�kv&�a�ɑ���-
��~��6��C�
��L���O�Y������,>�Вzo%����G�j���Zz����rn��ï�>K?�,M|�^�����僙خ+���HYM�X�e�O�5R���}1�>PA�{�\I�wB��8̺0���ɕ(_�:'�}3J�˖jX[���F���s1�=Er'���i͵�Z[8�y���?�L��D�t7v���m �?�����t�C��d����� c�2hA���+����H��LgӘ{���EȖg[�`=���^��t���m��g]��um},ȼ ����7::-.��鸳!}Y;��l �o���~Ӹ�c<⽚�F��#���M�z��p��uX @xo�=�	Bnq�����$�u�oo_Z���!	IE�H���M�Ldt�aY���qL;Rg�����Z�`�'��Xey/���/4�L�h�v����I`e�mC�(��F�QL�����h�?���#��>��szJ�נ7���Kϴ`5�Vo��U�,�������%"�^� �݌5A<�`��w��97yuY��b,u�c��O��Of78�����}�Wr��wz�8zF+�_s��J�<�Z��T|�ߢ��t	q%�SSE���
*ȗH��V�T�]��	I���dc�vt�K��z�)o9@�����躠����dl٪��0�s=_�pZ�)6��U�KѼn����u��&=/����w��s-������a�����ڳp��JJ�FO�b��9^�Mm�����������c<H0���U|i-w��i%vM�V��ڧ]_ʈ���$r�i��'�Z�;���<��d�e�g��<����O�ypA���b��Dº�ؐB��S�}T��fl�����3Q<\7��F���oJ�MO3U~�XƜ�#����CgT�	h�lNO�09NN��[ޭ�6]�̱��uc�������H��,/Kg�r����d>�DUqf���-(c�������?H��?��������4�4u&��Ē�(~���6@gwN����ꎐ�^)?ju��m-%tk��C�5��|�/@�����A݈��B�g�ϲ�a����@}����B��� H��;��9�Y-�W B�#�ɪ�]SOۈ��\�h�l���Ƕ6)�t0�����`� 8Ŏo�@R;�/t��&�N<!:�<�	ZN�܅�������I>n��5�҇������:��?�Խ;�揯�U�/uE]�����D?⭷ ?_�I����r8w���^�8g{'�e���8Ԫ����#�O���/Ux�IU�	t�KECFE �kc�I���#������G��D2}G�%�Y�UF��~=����u�l�]�]W3٬��y�J�ZGF��^Z�K�0|Z9!�^���Ǳ�"o�e�jsJ����k,e�Y�
ig�q�>;980ķ�8Zd��a�0=�=j+���t����ԭ�:$�*�Xȶ!�f�;�-�@0x~��?Ow\~^��
�t�l�㕅�Ԃ-����L�PW��#FE�}����A1~4w����y� ��! ��r�Pźs!"��m���>P���:_���	G� ����)+�}+Q	� �+G���{!��c���L3��y���1(�X���!'+�M�۰�`1y�LXx����k;擹�	B��T������Y�	��H��=�����-.w�ãذ����~��>h�S���LEWCj,�������hv�d5�1H� G��
��>7�G$�+�D��,���H�5ղB]�����l:pL���(��;y��� ���e�t�]%��}'!) ��h$�SN�\��#��ĸ?���,��7O��qjs�y�L�A�9��Jn87[��n+M�?���9oU{�RR[���ЇF5H[�tF������*U sb	`'��L�׻�ǛC�,�N�0ԡO�_I�.ͭ��lR��@�q�U�u�ExQ�_��6�\A=>��i*4�����8��%;�8�= ��Ѥ�o]8w��/��&V-�|ww
���n �o��Ž������@�����Q����8��v��Y�QM����������䲅�W�w�~)aH��Pœ����f8����zl�;Β�BU�NۤÚf�gԖ�g߹dv.����7�I6�z�ސ�	ԟ_���������X�ޘz� ���K>�䳀Po�l�x�d8'�Rwa������wj�Ay����}���S�s(_�t����#�ގ'e��*G�X0��Rn�nD��r�W�>e���g�9�WI���G�o��s��@�>r�cO�]I��`;�!8�bKACL\*�e�q.����0��wx�����_;�/�̘V�
�MB�}���P���`��F�&�_����;v�f�s_w�Sfi�3�T.lA�W,���y3�'�9D��%����,�!m�܃�M�2[n�i&�
P!�sG;��c��ބ��e��i����Ay��������43�Ex�Fի;I ؖMA�4�����O!W��X^.c�P/���'E�3�t�3C�ɲ7c��E��x����
G��J���5f�\�L}� �̔zgu�K�۳8����8�Yz�����ސ��S���@���5�^��7�d��p�^�����ܘ�Fa���bp��Ԩ��]	�x�(�J�VФ�QкD��z}аB�P"�Ȣq�V��*�8�&36ڠ��2g�!�y����t�E(�[��=	NVFޥZ��h-Nqc��C$����!�ĺχ�f__*�Կͧ�_n	��Ó�}C�Z�5��
jX֨@G�?���lV<ix��>��Wn���Ԣ��	�̌��T��Ga�}�~֔�[�2��^����׵����u+���
_������Z�n5Oa13[�4o��\�#3-�p^�Sxu�r> �J�u݃֓�QU�7�vpQ��^(Y�� L�v�,�lLJO<�h����Iz;�؀W_� ��zo�c�*��(���K4���n��j^T>v��W-o5b �G��-�d�	�������������6��.ʔ@��I�$�Q���f�gX9���v�K�����@:UBY�� �L���GXt[�63��j�'��9=7\��T;�` �.ph2Exym���1���wd�3~�Dd>Epv�[��D"����%E�L����*r���K��b�Ҧ�L����+�L�g�a*�1�iRp+
���y�a�8����Y������|⹭4f���֪Xa��x%����+EC���Ig�hwб��9�(�{Wca�V����h�����]�:A{�ۛ@�c��	����]j�C�e4��(>��j_�"w]����E�m�����f��N���i�E�M����r�K�.�RMu.����h��F�����)�Y-���%��ȰKw4�~PE�`˚��N o ��J���qbY��(Lr�����v�K��~��6�y�Nc#��.j�	���~& ��jqb��.��!o)	L�;W��x�=�ɕ�� �?���#����M|���.��g��"�.%�Ϝ�EL��e��|)����隝���:s��鈻0"N=gI'_�\(�g�܆�?֊�� Lhtm�~[a��ޏ�?�HF=n�����i�y9H']��/\
�8���,�t8a�E�#U؍at��7�)݊��s�Xn�1��ue���]���w=� �
j�����<��	�[��g�+H���������dRv~b�3 �V~*p�Oj
&��b���>F!���;�O33����@^�+����q��T��F8s7��ʉ�	���T�jV�i�J��H	Z�Z�G��ȅ7L�E�2�+2��q��|������l����yWj$n��~��\��F��+\����cZ�3>^WFf:P^*��[�����A��~ �Ҽ�4��_����8�����4�>6��Ꮻ"���{@,�ȑ�/I"�[]�=�����	F��}�F�^�\������O�A�N˂u�F�#����I1�AD�Ka��������h�2慴��Xq��M��C����y����$�����L�M��cor�b�5_sAy���m�ucՏG�ʵ���$&V��nvw��W���-����1�I�Ցof�/�sF�B����@|1Y�Z\��*q�hߎ�s#�2欔���ت4RW:DG�:
0)������j����K��c�2m]�a{�G�������!Ej�MtRڮ�V�AC�|d��+��ǝ����jy-�A�!M��#������i��\|Nz�u8-I^�5_к5��,��XP|�DŢ�,P�th�\eL-kW�����<��K�.א`3��c4�R?�a�0�.i���J�^f�sy=�� ��;|�pyR߿�YXr���b��	e�LS;}�>%R�[�X����-+�~t��E15'����a�V�������=!����f���:�"f+�2��ι�6)�-oX6�d2�
Ļ�׺�|�v-���i����~e�7�رț�n�*��H}w��Om�հ@��F��
ʈ&�>K�xl�+�4�;M��ڜK �j5����m���ᶜ(;����K��5�g�y��z�e����MuF �M���L��N)���i��0���t�)��A��<����oE�ZD3�5x69[S2�
�x��&���wO6�8�)�e��,�4q�bx)�Ni2�)�����N&��*X������*T f�I�XP�V�־�:IwR�du�:(�wV!�G����v����֜�3�3�V�DÉ�XU4J.1�.�{)~�.*�u��?�x��X?�n�C?n�ro�Y����Ʃ(��J�Y�)��U�׭�t���%%�M2�~o�Pwh7:���N6U���g���WT����t8+�X.���%�;M�/^�=ή����C��#�&���!���M�ƃ�i<٢��aJ4�]���i�Y)˙HDn!3�,�j�À�q�p{�ԁ16f�i�����%6'S���h2��*G�2b*id}Yn-���&z�dp�����tBU!���V��"m����� ;�������(�٭+����8,|Rt����Ȁ��x��f~�4���x�=��ȳ��d��[E.��o�hC�c\��$��x���ӕԦ�S]�\�.�����G�}W$��E
�'�!�~���?"�%>���Ψ��s�2��l���.\�Oq
G�hCsd=O[Ĵ�p����@��{w�~��Se��_�!,K��� �.�� ��i9)�w�7JWk�P�n%��#)E�DT�-���*�
�Aן�B�	l�����)m�Е�vA�������#��adIhK!(|d���1� ���>�JA��������z�ֺ	oC-2�ǥ�[��l"���H���m���E�0�n��ˬ�s���^�g}�!(e����6����3�N��դ)I��p;�@�"��G��f"8�s��G��q�D��\�[ם�!Ç�� �%'����+��dQ���ݬMl�����[>[e��[=�5�K>~y�)�L�	Y�(�=��l����߄f�(|�|6���u3ŧ�}p-�*j��f̭�k};u��:X��U��X߰��*|0,	'�O��-��Z�G�3^�w'+� �Ҧ��0�p	���K���D��_;-������qs��Hh�S�M	Ւ�����1̂���FP���ϟ��"}�B�>��zd�E�24�,�^�T����
q�_m-.o=�����/��bj[q%Dtm毣���B�\��#u	�b�=N��i�Iy��9�4S��3tEV+I�B�*ǮT'=9�d.W�dǗ��I��@~�9xV�b"�;�8��a�Yl���� T�AT& �΀"m�)
�F�	�f6{�Y^��:;�O�h(y�i��$q-w���L
ޟ��$�f(��,�g�_:� �q��g3?K��������f�3��9P���s���p�IL]�� }�𤋮��#�ly5=����fZ�.�����h�Q2���&ك/��!��KR2�H�h	L1d�}�'�@�e�AA���x3�B�<M���w&�.hJkT��/�π\�GI'Dk� ��=d&=۸d&%}	mRMƼdh��J��Y)7Jw@h�ߝs�5�
!��Y���A9��(#|J�N6FHq aJ�E�@ў�Y �ê��R�b��(�p�뻕��{N�>�O\O�R��Uu�'�#�Q�eH�`��+9�m���Y���I�#���-�K�v�U��+�
�_wuq ���g�DL(7��|���`��,Q��}�,�Bʆ�XY�c�R]�u�hu<ꕟpT7c��|�(P׫ѣA�%��zR��Ɂ�.�2G�������%��}�,g~�;�2<Ľ���4�J_W�� ����R��^�bK���J��g�ju��*��6+)��x�)�K�n�����WC6ց�����$8!ф����!����ai|ל�`��>�/�tNG��|&��L��Z�H�#��D��"g�P}�]6�q��CJ���׺�!�T�S��-`��9��\
ʽ$��C~	KAƉrI��T�لY�]���A�X�#��9b� ��գ���#.�sF�2�]6�r��	%^_��\م�3�Cu�Ir�A!�TÆ�r��:�}��$��g9�y<��w��Ì�'�L�'΢$JG�7�pdX�hY&�o�WP���)d�CW
U�N6�LϣԥFs��������Gx4%�V�K�p1iBzj$[R��a
�{�F�7!m'���J�p�{gN}�V����bP�4�댔��P�N�WZ[lfQ�#���UN2TrCrAs-@&_��/U`�[��{ț�j�z�S�[�~s!.�|y��v����#�k&�.ԫU���i><e�� �]����&��;U��Cژ�ZՈ#G��_��s2��*n���@\@f20o8�1g�z?a��oL�=)��Z�Ϛ�E$����Z	 dc�'��k�SKW��im� 5��z&Q>���Y��D-��'�l�ָD�.Z��4�!0�чo�	sD�)z�c��H&"X�U�8�2�����uR���B-F���F�����J�F��8;K�K���A,ﰇv��1'N���U�/����p��L/��a*N��~�p��"q�+��8U��tv�P�t����d}u�;<է'_�n��\1\���8��[���j�fѺ}L��I�1�§��7y��MK�z>��ʥBD��}��Cg��m��Á(�ӉYN�����f��_^;Ϝ�G.�t�-H�Q_�{<Ƀ��m�$"�/17��F�MϮ������Z���n��D�ҹڶ|�b��má�S�5�] �ႹK�K��(��C�l�.	�\n����~�oVYB��A�؁T`y;�,}˕Wܸ�-��Vp���W�2W!����<z�nm�0��kV�=;�t����h�B��4^����.%�1�{�L4����iCb܈cz�+G�|��n��1�fv�:���)d�J����������̥ƻ��|�����/��_����0���.�_������K������]#V��p9�s��d�П]Fr©���9�F@�>��
 #D��6��Xɲ�L��|$��B�M���c��q@�9h�k��q�B|^�����q0_x�ĀW�{$yEӡ:�tK��&�u?��r��{���a��hc&9~�7��V�Kh}w�ᄿw?b���$^,n�� �_��FTˡ��Wb���>�mU���{�4�v��0g�^�np'tU �MV�#;RO�g.�R	����u��*���ȶ S����bc%�F�5
\rD�ٳ���1?���W���⋬���B��(�XȎ$�s+hbF�����~�6�z+�P�(�V���V�M~yA�X&[T����-�jo+���=�yJ�d��"�I_|�X��D�)���`�
�!�A=AT!}e�(9�R�|��z� 
�wL�9��j<0O��9�Rw_�3�(��͹π�$���΄�ۣ�����U�!s��&��;���N�p{DQ{��T��Z�f:c��\] �@Ac���4�E�g��c�O�H�a�`��� �Ѕ�8ֈPO
FX]�՟��J*:[w���{��d�0ҕB���J��*y��)�p&J\�����A���2:d.�\!��j0 >�O󅄒J����9��Ț�7Ҋ@ع�56]�N@_�l�2or���gB�މ;�v����S|4m��(-��%�=$�Z�Á��'JаޗƌQ�0��h�����j��R#9�k���
)^f�GL�����oe�ȵ~����RŊ�J7Z�=�0]M�Y#]��W�V�\_"��+��ݒQ\V��cl{u����Y�$�Q�MyR��B-=�^�A�/����tF�m1�6uP!������e�Noeyd�T[$�&<�z*��ݟk8�᝸hQ���;[P���KlTsC�k2�>���br�f6�a��2� �<����\hؽ��m.;�� ^6���a���翞�N^��66T=cs�!F+��$ '����=��3�y�j��H��<���+�l$`V���a��d���~�W[^)�y�u�in�_�9��k�3������'���I;;Fh��ִ�6�	��VC�5_*7~؜L3�x��,	-�